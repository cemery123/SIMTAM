(* use_dsp48="no" *) (* use_dsp="no" *) module top #(parameter param290 = (7'h41)) (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h7e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire3;
  input wire [(5'h14):(1'h0)] wire2;
  input wire signed [(2'h3):(1'h0)] wire1;
  input wire signed [(3'h7):(1'h0)] wire0;
  wire [(5'h13):(1'h0)] wire289;
  wire signed [(3'h5):(1'h0)] wire288;
  wire signed [(5'h13):(1'h0)] wire286;
  wire signed [(2'h3):(1'h0)] wire12;
  wire signed [(4'h9):(1'h0)] wire11;
  wire [(2'h3):(1'h0)] wire10;
  wire [(3'h6):(1'h0)] wire9;
  wire [(4'hf):(1'h0)] wire8;
  wire [(5'h11):(1'h0)] wire7;
  wire signed [(4'h8):(1'h0)] wire6;
  wire signed [(5'h12):(1'h0)] wire5;
  wire signed [(2'h3):(1'h0)] wire4;
  assign y = {wire289,
                 wire288,
                 wire286,
                 wire12,
                 wire11,
                 wire10,
                 wire9,
                 wire8,
                 wire7,
                 wire6,
                 wire5,
                 wire4,
                 (1'h0)};
  assign wire4 = ((^~(~{wire0, (~&wire3)})) ?
                     (^~(($unsigned(wire1) | (wire0 ?
                         wire0 : (8'had))) | (8'ha7))) : (~$signed(wire1[(2'h2):(1'h0)])));
  assign wire5 = wire3[(4'h9):(3'h4)];
  assign wire6 = ($signed((wire1 ? $signed(wire2) : wire0[(1'h1):(1'h0)])) ?
                     (($signed((8'ha0)) & (8'haa)) >> $signed(wire5)) : wire5[(3'h5):(3'h4)]);
  assign wire7 = $signed($signed($signed((~^$signed((8'hb0))))));
  assign wire8 = (-{{((~&(8'hab)) ? (~^wire4) : (8'hb2))},
                     ({$unsigned(wire5)} ^~ (wire3[(1'h1):(1'h1)] ?
                         (~wire3) : (^wire1)))});
  assign wire9 = wire8[(3'h6):(2'h2)];
  assign wire10 = wire2;
  assign wire11 = ($unsigned(((^(wire8 ? (8'ha8) : wire8)) ?
                      wire4[(2'h3):(2'h2)] : (wire3[(4'h9):(1'h1)] ?
                          (wire7 ?
                              wire0 : wire10) : wire10))) - $unsigned((wire0[(3'h4):(1'h1)] >>> ($unsigned(wire8) ?
                      $unsigned(wire8) : (wire9 ? wire5 : wire0)))));
  assign wire12 = (wire0[(3'h4):(1'h1)] ?
                      wire2 : ($unsigned(($unsigned(wire7) <= wire9[(3'h4):(3'h4)])) >= $signed((|wire1[(1'h1):(1'h0)]))));
  module13 modinst287 (.y(wire286), .clk(clk), .wire16(wire5), .wire15(wire8), .wire14(wire2), .wire17(wire11));
  assign wire288 = $signed(wire1);
  assign wire289 = $signed(((^(~|$signed(wire11))) - ((~&(~|(8'h9d))) << ({wire4} ?
                       (-(8'hb1)) : $unsigned(wire288)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module13
#( parameter param285 = ({(^~(^(+(8'h9f)))), ((&((8'hb4) ? (8'ha9) : (8'hb8))) >= (!(8'had)))} ? ((((~&(8'hbf)) < {(7'h40)}) ? (8'hb7) : (&((8'hbf) ? (8'hba) : (8'hb8)))) < ((((8'hb5) ? (8'h9d) : (8'ha9)) >= ((8'hb8) ? (8'ha6) : (8'h9d))) >= (~(^~(8'ha7))))) : (({((7'h44) ? (8'ha0) : (8'hb2)), ((8'ha9) | (8'hbc))} ? (((8'haa) ? (8'hb4) : (8'hbd)) ? ((7'h43) || (7'h42)) : (|(8'ha6))) : (|{(8'hbc), (7'h43)})) ? ((((8'hae) ? (8'hb1) : (8'hb7)) ? ((8'hb4) ^ (8'hab)) : {(8'hbf)}) ? (+((8'ha4) ? (8'hb4) : (8'hae))) : ((^~(8'h9f)) * (8'haa))) : ((~|{(8'hb6), (8'hb8)}) - (&{(8'hb7), (8'h9c)})))) )
(y, clk, wire17, wire16, wire15, wire14);
  output wire [(32'h15e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire17;
  input wire [(5'h12):(1'h0)] wire16;
  input wire signed [(4'hf):(1'h0)] wire15;
  input wire [(5'h14):(1'h0)] wire14;
  wire [(5'h11):(1'h0)] wire284;
  wire [(4'hb):(1'h0)] wire283;
  wire [(4'h8):(1'h0)] wire281;
  wire [(4'ha):(1'h0)] wire206;
  wire signed [(3'h7):(1'h0)] wire205;
  wire signed [(3'h7):(1'h0)] wire204;
  wire signed [(4'hc):(1'h0)] wire203;
  wire [(4'hc):(1'h0)] wire202;
  wire [(4'he):(1'h0)] wire201;
  wire signed [(4'hf):(1'h0)] wire200;
  reg [(2'h2):(1'h0)] reg199 = (1'h0);
  reg signed [(4'he):(1'h0)] reg198 = (1'h0);
  reg [(4'hd):(1'h0)] reg197 = (1'h0);
  reg [(3'h6):(1'h0)] reg196 = (1'h0);
  wire [(3'h4):(1'h0)] wire70;
  wire signed [(5'h13):(1'h0)] wire29;
  wire signed [(4'hc):(1'h0)] wire28;
  reg signed [(2'h2):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg25 = (1'h0);
  reg [(5'h11):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg22 = (1'h0);
  reg [(4'h9):(1'h0)] reg21 = (1'h0);
  reg [(5'h11):(1'h0)] reg20 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg19 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg18 = (1'h0);
  wire [(4'hb):(1'h0)] wire72;
  wire [(4'h8):(1'h0)] wire104;
  wire signed [(2'h3):(1'h0)] wire194;
  assign y = {wire284,
                 wire283,
                 wire281,
                 wire206,
                 wire205,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 wire70,
                 wire29,
                 wire28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 wire72,
                 wire104,
                 wire194,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg18 <= {$unsigned((~((~|wire16) ? {wire14} : {wire16, wire16})))};
      if ((8'hbe))
        begin
          reg19 <= (~($unsigned(($unsigned((8'hba)) && reg18[(4'h9):(1'h1)])) * ((reg18 ?
              (wire17 ? (8'hba) : wire14) : $unsigned(wire14)) != ((wire17 ?
              reg18 : reg18) >= (!wire16)))));
        end
      else
        begin
          reg19 <= ((^~(((^wire14) ? (8'haa) : {wire14, wire15}) ?
              $signed(reg19) : $unsigned(wire17[(1'h0):(1'h0)]))) ~^ (~$unsigned((~^{(8'h9d),
              reg19}))));
          reg20 <= (7'h42);
        end
      if (reg20)
        begin
          if (wire15)
            begin
              reg21 <= wire17;
              reg22 <= ((&wire14) ?
                  (8'hb7) : ((((7'h42) ? (wire14 ? reg20 : wire14) : (^reg18)) ?
                          $signed($unsigned(reg21)) : (8'h9c)) ?
                      $signed((~&(reg20 ? reg19 : wire14))) : wire16));
              reg23 <= (8'had);
              reg24 <= (^~(~^$unsigned($signed((reg20 ? wire14 : reg20)))));
            end
          else
            begin
              reg21 <= {$signed($unsigned(reg21[(3'h6):(2'h3)]))};
              reg22 <= $unsigned(((wire15[(3'h4):(2'h3)] >> $unsigned($unsigned(reg20))) ?
                  $unsigned($unsigned((wire17 > reg22))) : (reg19[(3'h5):(3'h4)] ^ {(wire16 ?
                          reg21 : reg22),
                      wire17})));
              reg23 <= wire15;
              reg24 <= ((reg23[(5'h13):(4'he)] ?
                      (wire16 != ({wire14} ? (8'hbd) : wire16)) : reg23) ?
                  {(|($unsigned(wire17) ?
                          (reg18 ^~ reg24) : ((8'hb7) ?
                              wire17 : (8'hb8))))} : ($signed((~&$signed(reg21))) < $unsigned(wire17)));
            end
        end
      else
        begin
          reg21 <= reg22;
          if (wire15)
            begin
              reg22 <= (wire17 ~^ (wire17 ?
                  (^~$signed((+(8'had)))) : (~^reg23[(2'h2):(1'h1)])));
              reg23 <= wire17;
              reg24 <= wire17[(3'h5):(1'h1)];
              reg25 <= ((wire15 ?
                  ($unsigned(((8'hb5) ^ wire16)) * reg18) : reg23[(5'h14):(5'h11)]) && (reg22[(4'ha):(3'h7)] ^~ $signed(reg21)));
              reg26 <= wire14[(5'h14):(4'hf)];
            end
          else
            begin
              reg22 <= $unsigned(((8'hb7) ?
                  (((reg23 | (8'hb3)) || $signed(wire14)) ?
                      (~&$unsigned(reg23)) : (reg21 >> (&(8'ha4)))) : (&(reg19[(3'h4):(3'h4)] ?
                      $signed(reg24) : ((8'hb3) + reg24)))));
              reg23 <= ($unsigned($unsigned(((^reg24) + (reg20 ?
                      wire16 : wire16)))) ?
                  $unsigned((reg25 ?
                      reg20 : reg26[(2'h3):(2'h3)])) : reg23[(4'h8):(1'h1)]);
              reg24 <= (~&$signed($unsigned($unsigned(reg22))));
              reg25 <= ($unsigned((reg22[(3'h5):(2'h3)] ?
                      $unsigned(reg23) : $signed(reg20[(4'h8):(2'h3)]))) ?
                  reg20 : (-$signed($unsigned((~^reg18)))));
            end
        end
      reg27 <= {{$unsigned(reg23[(3'h4):(3'h4)])},
          ($unsigned((~|(reg21 ?
              reg26 : reg24))) * {$unsigned($unsigned(reg18)), wire16})};
    end
  assign wire28 = $signed({$unsigned(((~|reg21) ?
                          (reg23 ? reg24 : wire15) : reg26)),
                      $unsigned($signed(reg21[(1'h0):(1'h0)]))});
  assign wire29 = (reg21 ?
                      wire14[(2'h3):(1'h1)] : $unsigned((reg27[(1'h0):(1'h0)] * $unsigned(((8'hb5) ?
                          reg20 : wire17)))));
  module30 modinst71 (wire70, clk, reg22, reg19, reg20, reg18, wire15);
  assign wire72 = {reg20};
  module73 modinst105 (.wire77(reg20), .wire76(wire72), .clk(clk), .wire74(wire15), .y(wire104), .wire75(reg24));
  module106 modinst195 (wire194, clk, reg23, wire28, reg26, wire72, reg20);
  always
    @(posedge clk) begin
      reg196 <= {$signed(wire28[(3'h5):(3'h5)]),
          ($signed(wire15) > $unsigned(wire28[(3'h5):(1'h0)]))};
      reg197 <= reg19;
      reg198 <= reg22;
      reg199 <= ({wire14} ?
          ((({wire194, reg197} + {(8'hb4)}) >> wire28) ?
              {(reg19[(3'h6):(1'h1)] <<< (&reg21)),
                  ((+wire17) || wire15)} : reg20) : (-$signed({reg25})));
    end
  assign wire200 = wire104;
  assign wire201 = $signed($signed(wire16[(4'hc):(2'h3)]));
  assign wire202 = {$signed((&(!$unsigned(wire70))))};
  assign wire203 = reg196[(2'h3):(1'h0)];
  assign wire204 = reg199[(2'h2):(2'h2)];
  assign wire205 = reg22;
  assign wire206 = $unsigned((($signed($unsigned(reg18)) << wire202) ?
                       ((reg196[(1'h1):(1'h0)] ? wire14 : {reg23, reg196}) ?
                           ($signed((8'ha6)) ?
                               reg20[(2'h3):(2'h3)] : (wire194 ?
                                   (8'ha4) : reg27)) : $signed($signed((8'ha3)))) : (((reg196 ?
                           wire15 : wire202) * $unsigned(reg27)) ~^ $unsigned($signed(reg196)))));
  module207 modinst282 (.wire211(wire205), .wire208(reg21), .clk(clk), .wire210(wire15), .wire209(reg23), .y(wire281));
  assign wire283 = {(reg196 < (~|wire29[(4'h8):(3'h4)])),
                       $signed(({wire204} ~^ ($signed(wire194) ?
                           (wire104 ? reg197 : wire15) : $unsigned(reg199))))};
  assign wire284 = (^wire200[(3'h5):(2'h3)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module207  (y, clk, wire211, wire210, wire209, wire208);
  output wire [(32'h34a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire211;
  input wire [(2'h2):(1'h0)] wire210;
  input wire [(5'h12):(1'h0)] wire209;
  input wire signed [(4'h9):(1'h0)] wire208;
  wire signed [(3'h7):(1'h0)] wire280;
  wire [(4'h9):(1'h0)] wire279;
  wire signed [(3'h5):(1'h0)] wire278;
  reg [(5'h12):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg274 = (1'h0);
  reg [(4'h8):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg270 = (1'h0);
  reg [(4'hc):(1'h0)] reg269 = (1'h0);
  reg [(5'h14):(1'h0)] reg268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg267 = (1'h0);
  reg [(4'ha):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg263 = (1'h0);
  reg [(5'h12):(1'h0)] reg262 = (1'h0);
  reg [(4'hc):(1'h0)] reg261 = (1'h0);
  reg [(2'h2):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg258 = (1'h0);
  reg [(4'he):(1'h0)] reg257 = (1'h0);
  reg [(5'h12):(1'h0)] reg256 = (1'h0);
  reg [(3'h4):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg254 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire253;
  reg signed [(3'h7):(1'h0)] reg252 = (1'h0);
  reg [(4'hc):(1'h0)] reg251 = (1'h0);
  reg [(2'h3):(1'h0)] reg250 = (1'h0);
  reg [(4'hb):(1'h0)] reg249 = (1'h0);
  reg [(2'h3):(1'h0)] reg248 = (1'h0);
  reg [(4'ha):(1'h0)] reg247 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg245 = (1'h0);
  reg [(5'h13):(1'h0)] reg244 = (1'h0);
  reg [(4'hd):(1'h0)] reg243 = (1'h0);
  reg [(5'h15):(1'h0)] reg242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg239 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire238;
  reg signed [(4'he):(1'h0)] reg237 = (1'h0);
  reg [(3'h7):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(4'ha):(1'h0)] reg234 = (1'h0);
  reg signed [(4'he):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg232 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg231 = (1'h0);
  reg [(4'hb):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg229 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg227 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg226 = (1'h0);
  wire [(5'h12):(1'h0)] wire225;
  reg signed [(5'h10):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg220 = (1'h0);
  wire [(4'hb):(1'h0)] wire219;
  wire signed [(5'h10):(1'h0)] wire218;
  wire signed [(4'ha):(1'h0)] wire217;
  wire signed [(5'h12):(1'h0)] wire216;
  wire signed [(5'h14):(1'h0)] wire215;
  wire [(5'h13):(1'h0)] wire214;
  wire [(5'h10):(1'h0)] wire213;
  wire [(5'h13):(1'h0)] wire212;
  assign y = {wire280,
                 wire279,
                 wire278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 wire253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 wire238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 wire225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 wire219,
                 wire218,
                 wire217,
                 wire216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 (1'h0)};
  assign wire212 = (wire208 && ($unsigned($unsigned($signed((8'hb7)))) ?
                       (((^wire209) << (wire209 - wire211)) || $signed((^~wire209))) : $unsigned((((8'ha6) + wire211) <<< (wire208 >>> (8'hac))))));
  assign wire213 = $signed($unsigned(wire208));
  assign wire214 = $signed((~&wire211[(3'h5):(1'h1)]));
  assign wire215 = $unsigned(wire214[(4'hd):(3'h7)]);
  assign wire216 = {(~|($unsigned($unsigned((8'hb1))) == (wire215[(5'h14):(5'h11)] ^~ (~wire212)))),
                       $unsigned({({wire210} <= (wire214 <= wire214))})};
  assign wire217 = wire215;
  assign wire218 = ({wire209,
                       $signed($unsigned(((8'hab) == wire212)))} & wire209[(4'he):(4'h8)]);
  assign wire219 = (wire217[(1'h0):(1'h0)] + $signed({($unsigned(wire212) ?
                           wire216[(4'ha):(3'h4)] : $signed((8'ha5)))}));
  always
    @(posedge clk) begin
      reg220 <= (~&wire208);
      reg221 <= wire208[(3'h4):(2'h2)];
      reg222 <= wire217[(3'h4):(3'h4)];
      reg223 <= (wire208 <= wire216[(4'h9):(2'h3)]);
      reg224 <= (wire214[(3'h7):(2'h2)] < (8'ha9));
    end
  assign wire225 = ($signed({($unsigned(wire213) ?
                           wire212 : wire213[(5'h10):(3'h4)]),
                       wire217}) | wire209);
  always
    @(posedge clk) begin
      if ($signed($signed((8'ha2))))
        begin
          reg226 <= $unsigned(wire216[(4'he):(4'hb)]);
        end
      else
        begin
          reg226 <= (^~(wire212 ?
              wire217 : ($signed({reg224, wire219}) ?
                  {(wire208 ? wire209 : wire217), wire214} : {(|wire208)})));
          reg227 <= (((~&$signed($signed(wire214))) ?
              $unsigned((!(wire213 ?
                  (8'h9e) : wire209))) : $signed(wire210[(1'h0):(1'h0)])) + (reg223[(2'h2):(1'h1)] ?
              (~^(~&wire219)) : (((~^reg226) ^~ {(8'hb4)}) < wire208[(4'h9):(2'h3)])));
          if (reg224)
            begin
              reg228 <= (~|(+((|{reg226}) ?
                  (wire215[(4'ha):(3'h4)] && (wire219 << reg221)) : (reg226[(2'h3):(1'h1)] != $signed((8'ha2))))));
              reg229 <= wire219[(3'h4):(3'h4)];
            end
          else
            begin
              reg228 <= ($signed(((~|wire217[(2'h2):(1'h0)]) ?
                  ($unsigned((8'ha8)) ?
                      reg224 : $unsigned(reg224)) : $unsigned((8'h9c)))) > reg221[(3'h5):(3'h4)]);
              reg229 <= reg228;
              reg230 <= reg228[(1'h0):(1'h0)];
            end
        end
      if (({$unsigned((wire212 - $unsigned(reg227))),
          $signed(((wire219 ? reg228 : wire217) ?
              (^~wire213) : (wire213 || reg229)))} != (reg221[(4'hc):(2'h3)] ?
          $signed((~(wire208 == reg226))) : ({reg223[(3'h5):(3'h4)],
                  $signed(wire214)} ?
              (~|{wire213}) : ($unsigned(reg230) < (wire217 ?
                  reg221 : reg229))))))
        begin
          reg231 <= (($signed(((wire219 ?
                  wire216 : wire217) != reg226[(3'h4):(2'h3)])) * (((wire225 ?
                          reg220 : reg226) ?
                      $unsigned((8'ha9)) : (8'haa)) ?
                  {(wire210 < wire225),
                      (wire214 ? wire216 : wire225)} : (~&(-wire215)))) ?
              ({((reg229 ? wire225 : wire213) ?
                      {reg220,
                          reg226} : (~&wire212))} | ((~|$unsigned(reg228)) ^~ reg220[(1'h1):(1'h1)])) : reg230);
          reg232 <= ((reg227[(4'hc):(4'ha)] ?
              wire212 : $signed(wire212[(5'h12):(4'hb)])) * {reg223,
              ($signed((wire208 > reg222)) || $unsigned(reg224))});
          if ((&(&((wire210[(1'h1):(1'h0)] ^~ (|wire212)) ?
              (!reg220) : reg227))))
            begin
              reg233 <= $signed({(reg230[(3'h6):(3'h6)] ?
                      (^~(reg229 == wire213)) : {(^~reg223)})});
              reg234 <= $signed(($signed(reg232) ?
                  reg227 : ($unsigned(reg228) * {{wire214, wire219},
                      (wire216 < (7'h43))})));
              reg235 <= $signed(wire225);
              reg236 <= reg233[(4'hb):(3'h7)];
              reg237 <= reg227;
            end
          else
            begin
              reg233 <= $unsigned(wire211[(1'h0):(1'h0)]);
              reg234 <= wire209;
              reg235 <= {($signed($unsigned((reg221 ?
                      wire214 : reg231))) < (($signed((8'h9c)) ?
                      $signed((8'ha5)) : $signed(reg222)) < $signed((reg237 ?
                      (8'hb6) : wire209)))),
                  ((~|$signed({wire215})) ?
                      (-((reg229 ? reg230 : reg222) ?
                          reg236[(1'h0):(1'h0)] : reg233)) : (&(~$signed(reg223))))};
            end
        end
      else
        begin
          reg231 <= $signed(wire208);
        end
    end
  assign wire238 = reg227;
  always
    @(posedge clk) begin
      if ((~|reg222[(4'hb):(3'h7)]))
        begin
          reg239 <= reg234;
        end
      else
        begin
          reg239 <= reg221[(4'ha):(3'h4)];
          if (reg231)
            begin
              reg240 <= (($unsigned(reg237[(4'hc):(4'h9)]) == ((wire225[(4'hf):(4'hb)] ?
                          $signed(reg235) : $unsigned((8'hbe))) ?
                      reg223 : {wire208[(3'h5):(2'h2)], $unsigned(reg227)})) ?
                  (~^{((^wire209) ?
                          (~reg222) : $unsigned((8'h9d)))}) : ({wire218,
                          reg224[(2'h2):(2'h2)]} ?
                      $signed(reg233[(2'h2):(1'h1)]) : $signed($signed($signed(wire219)))));
              reg241 <= (^((((reg240 ?
                      wire225 : reg222) <= wire238[(1'h0):(1'h0)]) * ((wire212 >> (8'hb2)) ?
                      wire215 : (wire209 ? reg236 : reg234))) ?
                  reg231[(3'h5):(2'h2)] : ($unsigned((wire218 && (8'hb3))) ?
                      (+(reg221 ? reg220 : wire238)) : $unsigned((~|reg240)))));
              reg242 <= {wire219[(2'h2):(1'h0)], wire208[(3'h4):(2'h3)]};
              reg243 <= reg223;
            end
          else
            begin
              reg240 <= reg232[(1'h0):(1'h0)];
              reg241 <= $unsigned(wire215[(4'ha):(2'h2)]);
            end
          reg244 <= {wire210,
              ((wire210 < $unsigned($signed(wire218))) ?
                  $signed({(~reg230)}) : $unsigned(reg235[(1'h0):(1'h0)]))};
          reg245 <= ($signed((reg237[(3'h4):(3'h4)] ?
              {reg239[(1'h0):(1'h0)],
                  $signed(reg237)} : $unsigned(reg226))) & $signed((+$unsigned(wire238))));
          reg246 <= (({$signed($signed((7'h40))),
                  (reg236 ? (wire225 <= reg221) : (reg233 ^ reg230))} ?
              $signed($unsigned(wire218[(3'h6):(2'h3)])) : $unsigned(($unsigned((8'hb1)) == $unsigned(wire217)))) & {wire217[(2'h2):(1'h1)],
              reg245[(5'h13):(3'h5)]});
        end
      reg247 <= wire208;
    end
  always
    @(posedge clk) begin
      reg248 <= wire210;
      reg249 <= wire215[(4'ha):(1'h1)];
      reg250 <= reg246[(2'h2):(1'h1)];
      reg251 <= (-$signed($signed({$signed(reg227), $signed((8'ha4))})));
      reg252 <= $unsigned(((($signed(wire212) != (reg229 ? (8'ha5) : reg241)) ?
          (reg233[(3'h7):(3'h7)] ?
              (reg244 >> reg227) : (reg233 > reg233)) : (&reg224)) ^~ $signed(($signed(reg222) ?
          (reg221 == wire210) : $unsigned(wire225)))));
    end
  assign wire253 = ($signed(((wire210[(1'h0):(1'h0)] ?
                           reg243[(1'h1):(1'h0)] : reg230) ?
                       (8'hab) : $signed({wire238}))) <= reg229[(3'h6):(1'h0)]);
  always
    @(posedge clk) begin
      if (reg229[(4'hc):(1'h1)])
        begin
          reg254 <= $signed($signed(((reg220[(2'h3):(2'h2)] ?
                  (!reg242) : (-reg250)) ?
              ($unsigned(reg223) ?
                  (wire253 * reg236) : reg242) : (|(~|reg221)))));
          reg255 <= (reg239 * reg236[(3'h7):(2'h2)]);
          reg256 <= (|reg250);
          reg257 <= ((~&(~&$signed($signed(reg227)))) ?
              reg231 : reg220[(4'ha):(3'h7)]);
        end
      else
        begin
          reg254 <= reg243[(4'hc):(2'h2)];
          reg255 <= reg242[(4'hc):(3'h4)];
          reg256 <= $signed(((|({reg240, reg241} > reg248)) ?
              wire215[(4'hf):(3'h5)] : wire215[(4'hb):(3'h5)]));
          if (reg241)
            begin
              reg257 <= (wire218[(3'h4):(1'h0)] >>> $signed((!$unsigned((8'ha8)))));
              reg258 <= $unsigned(wire217);
            end
          else
            begin
              reg257 <= reg258[(1'h0):(1'h0)];
              reg258 <= reg242[(5'h15):(2'h2)];
              reg259 <= (((wire208[(3'h4):(3'h4)] + reg221) << ({wire214[(4'hf):(4'hb)]} ?
                      ((+wire215) ?
                          ((8'ha3) ?
                              (8'ha4) : wire208) : (wire215 - reg249)) : $signed(reg245[(1'h1):(1'h0)]))) ?
                  ((wire210 < reg230) ?
                      {(~(reg231 ? reg245 : reg220)),
                          ((reg233 ?
                              wire238 : reg222) >> (wire218 >> wire225))} : $signed(reg222[(5'h10):(4'hf)])) : reg243);
              reg260 <= reg254;
            end
          reg261 <= $signed($unsigned(reg224));
        end
      reg262 <= $unsigned(($unsigned(({reg247, reg255} > $unsigned(reg221))) ?
          {$unsigned((reg257 || (8'hb1)))} : (reg250 ?
              (reg257[(4'ha):(4'h8)] ^~ (!wire218)) : $unsigned((reg232 < reg250)))));
      reg263 <= (|(($unsigned((wire214 ~^ reg241)) ?
              ((wire218 ?
                  reg237 : (8'h9d)) <<< (reg243 < reg245)) : ((!(8'h9c)) ?
                  {reg222, reg256} : (!(8'hb6)))) ?
          reg241[(2'h3):(1'h1)] : $unsigned((~&reg222))));
      reg264 <= (reg258[(1'h0):(1'h0)] >= $unsigned(((wire218[(1'h0):(1'h0)] + reg259) == $unsigned(reg231[(2'h3):(2'h2)]))));
      if ($unsigned(wire214[(1'h1):(1'h1)]))
        begin
          reg265 <= (^(wire218[(4'hd):(2'h3)] ^~ $signed($unsigned((!reg241)))));
          if ($unsigned($unsigned(reg241)))
            begin
              reg266 <= (^~$signed((8'hb3)));
            end
          else
            begin
              reg266 <= $signed($signed((^~(wire225 << $signed(wire213)))));
              reg267 <= ((reg256[(4'h8):(1'h0)] ?
                  $signed($signed($signed(wire253))) : $unsigned((^reg260[(1'h0):(1'h0)]))) >= reg246);
            end
        end
      else
        begin
          reg265 <= reg229[(4'hb):(2'h2)];
          reg266 <= {$unsigned({$unsigned($signed((8'h9c))),
                  wire210[(2'h2):(1'h0)]})};
          reg267 <= (|$signed(wire213));
          reg268 <= (reg249[(4'ha):(3'h4)] <<< $signed($signed($unsigned($signed((8'hba))))));
        end
    end
  always
    @(posedge clk) begin
      if (($unsigned(((~&(8'hbf)) | wire209[(4'hb):(1'h1)])) ?
          {((!((8'h9f) ? reg245 : reg234)) & $unsigned((&reg259))),
              $signed(((reg223 <<< reg235) ?
                  (^~reg252) : (reg261 <<< wire210)))} : $unsigned((^(8'ha2)))))
        begin
          if (((reg234[(3'h7):(2'h3)] <<< $signed((reg239[(1'h0):(1'h0)] && reg233[(1'h1):(1'h0)]))) + $unsigned((wire219 ?
              wire212[(5'h11):(3'h6)] : ($unsigned(reg234) * $unsigned(reg243))))))
            begin
              reg269 <= {$signed(((reg252[(3'h6):(1'h0)] >= $signed(reg244)) - ((reg258 ?
                      reg248 : reg248) << {reg255}))),
                  (~^(reg267[(2'h3):(2'h2)] != reg243[(2'h3):(1'h1)]))};
              reg270 <= $unsigned($signed($unsigned(({reg248} <= $unsigned(reg268)))));
              reg271 <= ({(reg251[(2'h3):(1'h0)] >>> {reg248[(1'h0):(1'h0)]}),
                      ((8'hb0) ?
                          $unsigned({reg270,
                              reg229}) : (^reg243[(3'h4):(2'h3)]))} ?
                  (8'h9c) : (-$unsigned($unsigned(((8'ha3) | wire218)))));
            end
          else
            begin
              reg269 <= (((reg224[(4'hf):(4'he)] << wire209[(4'hb):(1'h1)]) <<< (8'had)) + (reg265[(4'h8):(3'h4)] ?
                  (8'ha0) : reg266[(4'ha):(2'h3)]));
              reg270 <= {(((reg239 - (~&reg250)) ?
                          ($signed((8'ha9)) >>> $signed(wire217)) : ($signed(reg237) < (&(8'hb4)))) ?
                      $unsigned(reg222[(5'h12):(4'h9)]) : ($unsigned($signed((8'ha4))) >>> reg267[(1'h1):(1'h1)]))};
              reg271 <= $signed($unsigned($signed(reg268)));
              reg272 <= reg251;
            end
          reg273 <= $unsigned((+(7'h42)));
          reg274 <= reg258[(2'h2):(1'h1)];
          reg275 <= $signed((((~^reg236) ?
                  reg251[(4'h9):(3'h4)] : $signed(wire216[(4'hc):(2'h3)])) ?
              ((reg263 + reg262[(2'h3):(2'h2)]) ?
                  (reg244 && reg227[(4'hd):(1'h0)]) : (^~(reg226 * reg233))) : $signed({(8'ha3),
                  (8'h9f)})));
        end
      else
        begin
          reg269 <= (reg234[(3'h5):(1'h1)] ? (!reg267) : (8'hba));
          reg270 <= {reg273, (~(^((~|reg245) <<< $signed(reg260))))};
          reg271 <= reg268[(3'h6):(3'h4)];
          reg272 <= wire212;
        end
      reg276 <= reg227[(4'ha):(3'h4)];
      reg277 <= ((-$unsigned(wire215[(5'h14):(4'he)])) ? wire238 : (8'h9d));
    end
  assign wire278 = wire218[(3'h7):(2'h2)];
  assign wire279 = (wire278[(2'h2):(2'h2)] ?
                       $unsigned($unsigned(reg251[(4'h9):(3'h4)])) : (8'hb4));
  assign wire280 = reg226;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module106
#( parameter param193 = ((~^{{((8'hb9) == (8'hb5)), (-(7'h44))}, ((-(8'hbd)) ^ ((8'hbf) ^~ (8'hbf)))}) < ((8'h9e) ? (((-(8'hb0)) >>> ((8'hac) == (8'hbe))) ^ {{(8'hbb)}, ((8'ha3) ? (7'h40) : (8'ha5))}) : (~|(-((8'hbd) ? (7'h41) : (7'h40)))))) )
(y, clk, wire111, wire110, wire109, wire108, wire107);
  output wire [(32'h325):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire111;
  input wire signed [(4'h8):(1'h0)] wire110;
  input wire signed [(5'h13):(1'h0)] wire109;
  input wire signed [(3'h6):(1'h0)] wire108;
  input wire signed [(4'hf):(1'h0)] wire107;
  wire [(4'hb):(1'h0)] wire192;
  wire signed [(4'hb):(1'h0)] wire191;
  wire signed [(4'hc):(1'h0)] wire190;
  wire [(4'h8):(1'h0)] wire189;
  wire signed [(4'he):(1'h0)] wire188;
  reg signed [(3'h6):(1'h0)] reg187 = (1'h0);
  reg [(4'hd):(1'h0)] reg186 = (1'h0);
  reg [(3'h6):(1'h0)] reg185 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg183 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire182;
  wire signed [(3'h7):(1'h0)] wire181;
  wire signed [(5'h12):(1'h0)] wire180;
  reg signed [(2'h2):(1'h0)] reg179 = (1'h0);
  reg [(3'h7):(1'h0)] reg178 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire177;
  reg [(2'h2):(1'h0)] reg176 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg175 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg174 = (1'h0);
  reg [(4'h9):(1'h0)] reg173 = (1'h0);
  reg [(5'h13):(1'h0)] reg172 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg169 = (1'h0);
  reg [(2'h3):(1'h0)] reg168 = (1'h0);
  reg [(4'ha):(1'h0)] reg167 = (1'h0);
  reg [(4'ha):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg164 = (1'h0);
  reg [(3'h6):(1'h0)] reg163 = (1'h0);
  reg [(3'h5):(1'h0)] reg162 = (1'h0);
  reg signed [(4'he):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg157 = (1'h0);
  reg [(2'h2):(1'h0)] reg156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg155 = (1'h0);
  reg [(4'ha):(1'h0)] reg154 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg153 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg152 = (1'h0);
  reg [(5'h11):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg150 = (1'h0);
  reg [(3'h4):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg148 = (1'h0);
  reg [(4'ha):(1'h0)] reg147 = (1'h0);
  reg [(5'h15):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg [(5'h11):(1'h0)] reg144 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire143;
  wire [(3'h4):(1'h0)] wire142;
  reg [(4'h9):(1'h0)] reg141 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg140 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg139 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg136 = (1'h0);
  reg [(5'h14):(1'h0)] reg135 = (1'h0);
  reg [(5'h10):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg133 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg132 = (1'h0);
  reg [(2'h2):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg129 = (1'h0);
  reg signed [(4'he):(1'h0)] reg128 = (1'h0);
  reg [(5'h14):(1'h0)] reg127 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg126 = (1'h0);
  reg [(5'h12):(1'h0)] reg125 = (1'h0);
  reg [(2'h3):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg123 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire122;
  reg signed [(4'h8):(1'h0)] reg121 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg120 = (1'h0);
  reg [(3'h6):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg118 = (1'h0);
  reg [(3'h4):(1'h0)] reg117 = (1'h0);
  reg [(3'h6):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg115 = (1'h0);
  reg [(4'hf):(1'h0)] reg114 = (1'h0);
  reg [(4'ha):(1'h0)] reg113 = (1'h0);
  reg signed [(4'he):(1'h0)] reg112 = (1'h0);
  assign y = {wire192,
                 wire191,
                 wire190,
                 wire189,
                 wire188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 wire182,
                 wire181,
                 wire180,
                 reg179,
                 reg178,
                 wire177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 wire143,
                 wire142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 wire122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg112 <= $unsigned(wire111[(3'h7):(2'h3)]);
      reg113 <= $signed($signed((~^((wire107 >= (8'h9f)) >>> $signed(reg112)))));
      reg114 <= (wire110[(4'h8):(1'h1)] ?
          ((^~(-wire108[(2'h2):(1'h1)])) * $unsigned(wire107)) : (|($unsigned(reg113) ?
              (-wire108[(2'h3):(1'h0)]) : wire108[(2'h3):(2'h2)])));
      if ($unsigned(wire109))
        begin
          reg115 <= (wire109 <= $unsigned(reg114));
          if ($unsigned($unsigned(reg115)))
            begin
              reg116 <= (^~reg113[(2'h3):(1'h0)]);
              reg117 <= wire110;
              reg118 <= $unsigned((($signed((+(8'h9c))) ?
                      ($unsigned((8'ha8)) < reg116[(3'h5):(2'h3)]) : (7'h44)) ?
                  reg116[(2'h3):(2'h3)] : wire108[(2'h2):(2'h2)]));
              reg119 <= $unsigned((($unsigned((reg116 ?
                  reg113 : wire110)) > ({reg118, reg118} ?
                  (wire109 ?
                      reg117 : (8'hb0)) : $unsigned(wire109))) - {(~|{reg112}),
                  ((wire110 ? reg118 : reg114) >>> (wire110 & wire108))}));
              reg120 <= $signed($unsigned(($signed(reg118[(4'h9):(2'h2)]) - (wire110 + $signed(reg112)))));
            end
          else
            begin
              reg116 <= (^~(($signed($signed(reg115)) ?
                      ((~|reg113) ? (reg113 ^ reg112) : reg120) : ((wire110 ?
                              wire107 : reg118) ?
                          (reg112 | wire109) : wire109)) ?
                  reg112 : $signed(((reg117 ? (8'ha5) : wire110) ?
                      wire109 : (~|reg115)))));
              reg117 <= ((($unsigned((wire107 <= reg114)) ?
                  ((reg117 ? wire111 : wire108) ?
                      $unsigned((8'ha4)) : wire108) : reg115[(4'hc):(1'h1)]) + (8'hb3)) > ((~$signed(wire109[(4'hf):(4'hb)])) - reg112));
              reg118 <= (({(^~$signed(reg120)), ((8'hb7) << (~^(8'hbb)))} ?
                      $signed(wire111) : reg112[(3'h5):(2'h3)]) ?
                  reg117 : ((7'h43) ?
                      ($signed({reg112}) ?
                          reg115[(3'h5):(2'h3)] : $signed((wire108 ?
                              reg113 : wire111))) : (wire110 <= ($signed(wire107) == reg112[(3'h7):(2'h2)]))));
            end
          reg121 <= wire111[(3'h7):(1'h1)];
        end
      else
        begin
          reg115 <= wire108[(1'h1):(1'h0)];
          reg116 <= wire108[(1'h0):(1'h0)];
          reg117 <= (+((^~reg114[(4'hb):(4'hb)]) + $unsigned(((8'hbe) ?
              $signed(reg113) : reg114))));
        end
    end
  assign wire122 = $signed(reg121[(3'h4):(3'h4)]);
  always
    @(posedge clk) begin
      reg123 <= {({{wire110[(3'h5):(3'h4)]}, (&$unsigned(reg118))} ?
              wire108[(1'h1):(1'h1)] : (|wire122)),
          reg115[(3'h5):(2'h3)]};
      if ($unsigned(((reg121[(1'h1):(1'h0)] ~^ $unsigned(reg112[(3'h5):(3'h5)])) ?
          (wire107[(4'h8):(4'h8)] ?
              (~^{reg120}) : {$unsigned((8'hb4)),
                  (wire109 ? reg119 : reg115)}) : $unsigned(((~^reg113) ?
              $signed((8'haf)) : wire108[(1'h0):(1'h0)])))))
        begin
          reg124 <= reg123[(2'h3):(2'h2)];
          reg125 <= wire108;
          reg126 <= ((^~wire108) ?
              $signed((8'hae)) : (|(({reg113} * $unsigned(reg119)) ^ $signed((~reg113)))));
        end
      else
        begin
          reg124 <= reg119[(3'h6):(2'h2)];
          if ({(~$signed($unsigned((^wire111))))})
            begin
              reg125 <= reg117[(2'h3):(2'h2)];
            end
          else
            begin
              reg125 <= $signed(wire109);
              reg126 <= (reg119[(1'h1):(1'h0)] ?
                  (8'had) : $signed($signed(wire107)));
              reg127 <= (^~reg114);
              reg128 <= ((~&reg114[(4'hb):(4'h8)]) > $unsigned(wire111));
            end
          reg129 <= (^(8'ha3));
          reg130 <= (~|$signed((reg114 - $signed($unsigned(reg115)))));
          reg131 <= reg116[(2'h3):(1'h1)];
        end
      reg132 <= (((reg124 * {wire111[(3'h7):(3'h7)],
              $signed(reg123)}) == (reg115 != $signed(reg118))) ?
          (reg123 ^~ (8'hab)) : $unsigned((&$signed($signed(reg121)))));
      reg133 <= reg130;
    end
  always
    @(posedge clk) begin
      if (({wire108,
          ($signed((reg115 ?
              wire122 : reg115)) <= reg121[(4'h8):(3'h5)])} != (8'hbb)))
        begin
          reg134 <= reg126[(3'h6):(3'h4)];
          reg135 <= reg114;
        end
      else
        begin
          reg134 <= $unsigned(wire108[(3'h4):(1'h0)]);
          if (reg133[(3'h5):(3'h5)])
            begin
              reg135 <= $signed((-$signed({$signed(reg119)})));
              reg136 <= ($unsigned(reg129) ?
                  ($signed(reg125) > (8'ha5)) : reg114[(2'h3):(1'h0)]);
              reg137 <= ((reg129[(5'h10):(3'h7)] << ((reg118[(3'h4):(1'h1)] ?
                  reg112[(3'h4):(2'h3)] : reg127) >= $unsigned(reg118))) > (^$signed(reg134[(4'hc):(3'h7)])));
              reg138 <= reg119[(1'h0):(1'h0)];
            end
          else
            begin
              reg135 <= (8'hb8);
            end
          reg139 <= $signed(((reg119[(3'h5):(2'h2)] & {(reg125 ?
                  (8'h9f) : (8'hb0))}) * {(^reg115)}));
          reg140 <= {$signed(((&$signed(reg121)) ?
                  reg126 : {reg139[(4'h8):(1'h1)]}))};
        end
      reg141 <= $unsigned(reg116);
    end
  assign wire142 = reg127[(5'h14):(4'h8)];
  assign wire143 = reg134[(4'he):(2'h2)];
  always
    @(posedge clk) begin
      if ({(reg116[(1'h0):(1'h0)] ?
              (^~reg120[(2'h3):(1'h1)]) : {reg114[(4'h8):(3'h4)],
                  reg124[(2'h3):(2'h2)]})})
        begin
          reg144 <= ($unsigned(($signed((reg138 ? wire110 : (8'hb1))) ?
              (~|{reg115}) : reg118[(1'h1):(1'h1)])) ~^ (reg137[(2'h2):(2'h2)] >>> wire110));
          reg145 <= $signed(((!(8'haa)) ?
              $signed({(|(7'h40)), $signed(wire142)}) : $signed(reg137)));
          reg146 <= (~^reg133);
          if (reg116[(3'h4):(3'h4)])
            begin
              reg147 <= (wire111 ?
                  (+(((wire110 ? reg134 : reg119) ^ (reg120 <= wire107)) ?
                      $signed($signed(reg144)) : reg128)) : reg136[(3'h4):(3'h4)]);
              reg148 <= (($signed(((~^reg140) ?
                  reg117[(2'h3):(2'h3)] : (~reg112))) + {(reg129 ?
                      reg129 : reg121),
                  ((8'hb6) ?
                      (7'h42) : reg145)}) + ((!reg121[(1'h1):(1'h0)]) > $signed(((!reg123) ?
                  reg120[(1'h1):(1'h1)] : {reg119, reg115}))));
              reg149 <= $unsigned((reg120 <= reg112));
            end
          else
            begin
              reg147 <= reg148[(1'h1):(1'h1)];
            end
        end
      else
        begin
          reg144 <= $unsigned($signed(reg114[(2'h3):(1'h0)]));
          if (($unsigned(($unsigned((|reg129)) || ($unsigned((8'hba)) ?
                  $signed((8'hbf)) : (8'hb4)))) ?
              (reg121 ?
                  ($signed((+reg129)) <<< ((reg145 ? reg130 : reg140) ?
                      (wire109 ?
                          (8'hb4) : reg116) : $signed(wire107))) : $signed({wire122[(4'h9):(4'h9)],
                      $signed(reg114)})) : ($signed((&reg127[(4'hc):(3'h7)])) ?
                  wire108 : wire122[(2'h3):(2'h2)])))
            begin
              reg145 <= reg134;
              reg146 <= $signed((-reg148));
              reg147 <= (wire122[(2'h2):(2'h2)] <= (reg126 == (reg136 <= $signed($signed(reg115)))));
              reg148 <= reg120;
              reg149 <= (8'hba);
            end
          else
            begin
              reg145 <= $unsigned(({$signed($signed(reg149)), $signed(reg127)} ?
                  $unsigned($signed(reg148)) : ($signed((-wire111)) ?
                      reg114 : reg146)));
              reg146 <= wire122;
            end
          reg150 <= reg145;
          reg151 <= $unsigned($unsigned(reg125[(2'h2):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      if ({(~reg132)})
        begin
          reg152 <= ({$signed(reg117[(2'h2):(1'h1)]),
              ($unsigned((^~reg116)) ?
                  reg144 : reg126[(3'h7):(2'h2)])} == reg141);
          reg153 <= ((^$unsigned((reg150[(3'h4):(2'h3)] ?
              $unsigned(reg132) : $signed(reg112)))) ^ $signed($unsigned($unsigned((~reg150)))));
          reg154 <= wire142;
          reg155 <= $unsigned(((~($signed(reg136) ?
                  $unsigned(reg151) : $unsigned(wire142))) ?
              reg121[(3'h4):(1'h1)] : reg133[(4'h8):(4'h8)]));
        end
      else
        begin
          reg152 <= {reg145[(2'h3):(1'h1)],
              (reg150 ?
                  (($signed((8'ha0)) ?
                      reg129 : (reg150 ?
                          wire108 : reg124)) <<< $unsigned($signed((8'haf)))) : reg127)};
          reg153 <= (reg121 ?
              ((reg141 >= $unsigned($unsigned((8'h9c)))) - (reg148 != {(reg114 ^ reg149),
                  $signed(wire122)})) : (!reg124[(2'h2):(2'h2)]));
          if ((^~(~|{(&(reg118 <<< reg114))})))
            begin
              reg154 <= (~^(({reg118[(4'ha):(3'h5)],
                          (reg154 ? (7'h43) : (8'ha0))} ?
                      ((~|(8'hbc)) ?
                          ((8'ha2) ?
                              reg153 : reg126) : (~^reg128)) : $signed($signed(wire122))) ?
                  reg133 : (reg133[(4'h8):(3'h6)] || (-(reg132 ?
                      reg119 : reg119)))));
              reg155 <= wire108;
              reg156 <= reg119;
            end
          else
            begin
              reg154 <= reg120;
              reg155 <= reg147[(2'h2):(1'h1)];
              reg156 <= {(8'hb4),
                  (!(((+wire109) ^ $signed(reg114)) > (8'ha9)))};
            end
          if (reg145)
            begin
              reg157 <= ((&reg121[(3'h5):(1'h1)]) ?
                  (((reg123 * (reg120 ? wire142 : reg146)) ?
                          $signed((reg154 >> wire143)) : reg145) ?
                      $signed($unsigned($unsigned(reg134))) : (($signed(reg115) != (8'ha7)) ?
                          (^~reg155) : $signed($unsigned((8'hac))))) : wire107[(4'hc):(3'h5)]);
              reg158 <= reg147;
              reg159 <= (~|reg157);
              reg160 <= $unsigned(reg153[(2'h3):(1'h1)]);
              reg161 <= reg129[(2'h2):(1'h1)];
            end
          else
            begin
              reg157 <= $signed($unsigned(reg161));
            end
          reg162 <= $signed((reg136 ?
              (reg158 > reg141) : reg138[(2'h2):(1'h0)]));
        end
      reg163 <= $unsigned($unsigned(({((8'hb2) ? reg127 : reg128), reg146} ?
          reg160 : {(|(8'hab))})));
      reg164 <= (($signed((reg128[(4'ha):(1'h1)] ?
              reg144[(4'he):(4'hc)] : (^reg149))) >>> $signed($unsigned((reg137 ?
              reg129 : reg113)))) ?
          $unsigned($signed(reg112[(4'he):(1'h0)])) : $unsigned($signed($unsigned((|reg159)))));
      reg165 <= (($unsigned($signed($signed((8'h9c)))) ?
          {(reg138 ?
                  (reg139 ? reg164 : reg154) : (reg153 >> reg164))} : {reg129,
              (reg126 < {(8'h9e), reg154})}) > (reg136[(3'h4):(2'h2)] ?
          ($signed(reg153) < reg126) : reg134[(4'hd):(4'h8)]));
    end
  always
    @(posedge clk) begin
      reg166 <= $unsigned(reg123);
      if ($signed(wire110[(3'h7):(2'h2)]))
        begin
          reg167 <= (($signed(($signed((8'h9c)) ? (~^reg124) : (~&wire110))) ?
              (^~({(7'h44), reg129} ?
                  reg153[(2'h2):(1'h1)] : (reg126 ?
                      wire111 : (7'h42)))) : ((reg124[(2'h2):(1'h1)] ?
                      (reg123 ? reg149 : reg123) : (reg154 ? reg134 : reg127)) ?
                  reg155[(4'hb):(4'h9)] : (reg145[(3'h7):(2'h3)] >> (+reg130)))) || (+(reg166[(3'h4):(3'h4)] == $signed(wire107[(2'h3):(2'h2)]))));
          reg168 <= wire143[(1'h1):(1'h1)];
        end
      else
        begin
          reg167 <= (+{$unsigned(reg116),
              ($signed($signed((7'h41))) != (reg120 & (reg126 != reg148)))});
          if ((-$unsigned(reg145)))
            begin
              reg168 <= wire111[(4'h9):(1'h1)];
              reg169 <= reg155;
              reg170 <= ((~|$signed($signed((reg121 ? reg126 : wire142)))) ?
                  reg168[(2'h2):(2'h2)] : (^{{((8'ha4) ^ wire142)}}));
              reg171 <= (reg131 ?
                  {($signed((-reg170)) ?
                          $signed({reg112,
                              reg133}) : reg168)} : $signed(($signed((8'haa)) ?
                      reg145[(1'h0):(1'h0)] : ((-(8'hb1)) ?
                          (^~wire108) : (^reg141)))));
              reg172 <= $signed($unsigned(reg167[(4'h9):(4'h8)]));
            end
          else
            begin
              reg168 <= ($signed($unsigned(($unsigned(reg164) <<< (reg147 << reg136)))) ?
                  ((reg135[(4'h9):(3'h6)] > ((reg150 ?
                          reg162 : reg152) ^ {reg169, (8'hb0)})) ?
                      reg155[(4'h9):(3'h6)] : reg116[(3'h4):(1'h0)]) : (~reg126[(3'h4):(3'h4)]));
              reg169 <= (wire122[(4'hb):(2'h2)] ?
                  {(8'h9d),
                      (reg120[(1'h0):(1'h0)] ?
                          (^$unsigned(reg118)) : $signed((reg114 < wire107)))} : $unsigned(reg151[(3'h4):(1'h1)]));
              reg170 <= $unsigned($signed({$unsigned((reg115 ?
                      reg113 : reg125)),
                  ((reg160 ~^ reg118) ? $unsigned(reg113) : $signed(reg172))}));
            end
          reg173 <= reg115[(2'h3):(2'h3)];
          reg174 <= $unsigned(wire111[(1'h1):(1'h1)]);
        end
      reg175 <= (+(reg114[(4'hc):(2'h3)] ?
          {($signed(reg137) == $unsigned(wire122))} : reg171[(4'ha):(4'h9)]));
      reg176 <= (((8'hb1) ?
          ($signed(reg136) ?
              ({wire110} <= $signed(reg164)) : reg113) : reg121[(2'h3):(2'h3)]) - $unsigned((&(((8'hb0) ?
              reg147 : reg114) ?
          $signed((8'h9d)) : $unsigned(reg163)))));
    end
  assign wire177 = (^~reg147);
  always
    @(posedge clk) begin
      reg178 <= (reg176[(1'h0):(1'h0)] ?
          (($unsigned(reg147) * $unsigned((reg112 && reg151))) ?
              reg130[(4'he):(4'he)] : ($unsigned({(8'hba)}) + reg137)) : reg156);
      reg179 <= reg155;
    end
  assign wire180 = (~^$unsigned({$unsigned($signed(reg165)),
                       {reg178[(3'h6):(3'h6)]}}));
  assign wire181 = $signed(((~(-(reg174 >>> reg165))) ?
                       ({reg178, wire143[(1'h1):(1'h1)]} ?
                           ((^reg126) > (~|reg176)) : reg149) : reg179));
  assign wire182 = ($unsigned($unsigned(reg160)) >>> reg131[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg183 <= reg166;
      if ($signed({reg134}))
        begin
          reg184 <= $unsigned($unsigned((((&reg150) ?
              (reg164 ?
                  wire181 : reg117) : (8'hb9)) <<< $signed((reg162 | reg114)))));
          reg185 <= $unsigned((((reg169 ? {reg174, reg178} : $signed(wire110)) ?
                  $unsigned($unsigned(reg176)) : (+$unsigned(reg175))) ?
              reg154[(3'h5):(2'h2)] : (reg116 ?
                  $signed($signed(reg153)) : $unsigned((reg127 > reg168)))));
        end
      else
        begin
          reg184 <= $unsigned((reg133 >= reg124));
          reg185 <= (reg165 ?
              $unsigned(reg179[(2'h2):(1'h0)]) : $unsigned((reg166 >> $signed($unsigned(reg127)))));
          reg186 <= wire109[(3'h5):(1'h1)];
          reg187 <= $unsigned({(8'hb4)});
        end
    end
  assign wire188 = (($signed(reg157[(1'h0):(1'h0)]) ?
                           $signed((reg157[(1'h1):(1'h1)] * reg172[(4'hc):(4'ha)])) : (^~$unsigned((+wire109)))) ?
                       $unsigned($unsigned($unsigned((~&reg175)))) : reg126[(4'h9):(2'h2)]);
  assign wire189 = (!reg128[(4'he):(4'hd)]);
  assign wire190 = (reg123 ^~ $signed($signed(reg139[(3'h5):(2'h2)])));
  assign wire191 = {$unsigned(reg153)};
  assign wire192 = $unsigned(reg140);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module73  (y, clk, wire77, wire76, wire75, wire74);
  output wire [(32'h12c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire77;
  input wire signed [(4'h8):(1'h0)] wire76;
  input wire signed [(5'h11):(1'h0)] wire75;
  input wire [(4'hf):(1'h0)] wire74;
  wire [(2'h3):(1'h0)] wire103;
  wire signed [(5'h14):(1'h0)] wire102;
  wire [(4'hf):(1'h0)] wire101;
  wire [(5'h13):(1'h0)] wire100;
  wire signed [(5'h15):(1'h0)] wire99;
  wire signed [(5'h15):(1'h0)] wire98;
  reg signed [(4'hb):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg96 = (1'h0);
  reg [(3'h6):(1'h0)] reg95 = (1'h0);
  reg [(4'h8):(1'h0)] reg94 = (1'h0);
  reg [(3'h4):(1'h0)] reg93 = (1'h0);
  wire [(3'h5):(1'h0)] wire92;
  wire signed [(3'h7):(1'h0)] wire91;
  wire signed [(5'h10):(1'h0)] wire90;
  wire signed [(4'hf):(1'h0)] wire89;
  wire signed [(5'h12):(1'h0)] wire88;
  reg signed [(3'h4):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] reg86 = (1'h0);
  reg [(5'h14):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg84 = (1'h0);
  reg [(3'h4):(1'h0)] reg83 = (1'h0);
  reg [(2'h3):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg81 = (1'h0);
  reg [(4'h8):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg79 = (1'h0);
  reg [(3'h5):(1'h0)] reg78 = (1'h0);
  assign y = {wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 wire92,
                 wire91,
                 wire90,
                 wire89,
                 wire88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire77)
        begin
          if (wire76[(3'h7):(3'h4)])
            begin
              reg78 <= $unsigned({$unsigned($unsigned(wire76)),
                  (($unsigned(wire75) && (wire77 ?
                      wire74 : wire76)) < (~&(wire77 >= wire76)))});
              reg79 <= ($signed(wire75[(4'hd):(4'h8)]) ?
                  ($signed((|wire75)) ?
                      reg78[(1'h1):(1'h0)] : (7'h42)) : $signed($unsigned(wire77)));
              reg80 <= {((({wire75, (8'h9d)} ~^ $signed(reg79)) ?
                      {(wire76 >>> reg79),
                          (-reg79)} : wire76) || ($signed(wire74) ~^ {(!(7'h44))}))};
              reg81 <= $unsigned($signed((+$unsigned($unsigned(wire76)))));
              reg82 <= $signed(($unsigned($unsigned(((8'hb6) ?
                      reg78 : wire74))) ?
                  reg81 : (+{(wire74 <= reg78)})));
            end
          else
            begin
              reg78 <= $signed((reg82 ?
                  {(!wire77[(2'h3):(2'h3)])} : reg80[(3'h7):(2'h3)]));
              reg79 <= $signed(($unsigned(((&reg79) ?
                  (|(8'haf)) : (reg81 << wire77))) ^ {wire75}));
            end
          reg83 <= $signed((reg81 | wire76));
        end
      else
        begin
          reg78 <= reg81;
          reg79 <= (^reg80);
          reg80 <= {(!$signed({$signed(wire75), (reg78 > reg80)}))};
          reg81 <= $unsigned(reg78);
          if ($signed(({wire74,
              ((reg79 & (8'ha7)) | (~^wire74))} << (!$unsigned(reg78)))))
            begin
              reg82 <= $signed($unsigned((reg78[(3'h5):(3'h5)] + $signed($signed((8'ha9))))));
              reg83 <= wire75;
              reg84 <= $signed((reg80[(3'h6):(3'h4)] ?
                  ((8'hbb) ?
                      $unsigned(wire77[(1'h0):(1'h0)]) : reg78[(2'h3):(2'h3)]) : reg78[(3'h5):(3'h4)]));
            end
          else
            begin
              reg82 <= {wire75[(5'h10):(1'h1)]};
              reg83 <= (wire77[(3'h4):(2'h2)] ^~ $unsigned((reg83 ?
                  (reg79[(4'hc):(3'h7)] ?
                      wire75 : (8'hb4)) : $signed($unsigned((7'h41))))));
              reg84 <= ($signed((~|{reg84[(1'h1):(1'h0)],
                  (~reg80)})) < reg80[(4'h8):(3'h4)]);
            end
        end
      reg85 <= $signed(({reg79} ?
          (wire74[(1'h0):(1'h0)] >> $signed(reg82[(1'h1):(1'h0)])) : {(reg81[(5'h11):(4'ha)] ?
                  ((8'hba) ? (8'hb3) : reg80) : (^~reg84))}));
      reg86 <= {$signed(reg79[(4'h8):(2'h2)]),
          $signed(($signed($unsigned(reg78)) < (^$signed((8'had)))))};
      reg87 <= {(-$unsigned({$signed(reg86), (reg81 ? reg83 : reg82)})),
          $unsigned($unsigned((~&{reg79, reg78})))};
    end
  assign wire88 = (~$signed({reg83, $unsigned((+reg78))}));
  assign wire89 = $signed((reg81 ?
                      $signed($signed((&reg79))) : (^(wire88 == $signed(reg85)))));
  assign wire90 = wire75[(1'h1):(1'h0)];
  assign wire91 = {(reg84[(3'h6):(1'h1)] ? wire89 : reg78)};
  assign wire92 = $unsigned((reg84 ?
                      ((+$signed(wire90)) >= $signed($signed(wire76))) : $unsigned($unsigned({wire77,
                          (8'hbd)}))));
  always
    @(posedge clk) begin
      reg93 <= (~|$unsigned((^$signed((wire76 && reg82)))));
      reg94 <= (8'hab);
      reg95 <= reg79;
      reg96 <= ($unsigned((((wire75 ? wire76 : reg78) & reg82) ?
          reg79[(4'hb):(4'ha)] : ((wire92 | reg79) ?
              $signed(reg80) : $signed(reg85)))) < (^(({reg86, reg82} ?
          wire91[(1'h0):(1'h0)] : (reg82 ?
              reg79 : wire88)) + (reg81 == $unsigned((8'h9c))))));
      reg97 <= {reg84, (~^$unsigned(reg95))};
    end
  assign wire98 = (~($signed({reg97, reg97}) ? reg85 : wire89[(3'h5):(1'h1)]));
  assign wire99 = ((wire89 && $unsigned(reg85)) ?
                      (reg83 ?
                          $unsigned($unsigned(reg86[(4'h8):(3'h4)])) : ($unsigned((reg81 ?
                              reg94 : reg84)) <= $signed($unsigned(reg85)))) : $signed((^(reg78 < (~reg87)))));
  assign wire100 = (wire75 & (reg81 & (^~reg85[(3'h4):(1'h0)])));
  assign wire101 = $unsigned(((|wire75[(4'ha):(1'h0)]) >> $unsigned(wire99)));
  assign wire102 = {($signed($signed(wire88)) >>> (-{{wire75}}))};
  assign wire103 = $unsigned(wire99);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module30
#( parameter param68 = ((-(({(8'h9d), (8'ha2)} == {(8'h9f)}) ? ((&(8'hb2)) <= (8'h9f)) : (+((7'h42) << (8'hb0))))) ? (~|{(8'hb5)}) : ({({(8'hbc), (8'haa)} >= ((7'h42) ~^ (8'hb3))), ((|(8'hae)) ? ((8'hb5) ? (8'hbb) : (8'hb0)) : ((8'hb3) ? (8'hb7) : (7'h40)))} ? (8'hb0) : (|{((8'hb9) ? (8'hac) : (7'h44))})))
, parameter param69 = param68 )
(y, clk, wire35, wire34, wire33, wire32, wire31);
  output wire [(32'h164):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire35;
  input wire signed [(3'h4):(1'h0)] wire34;
  input wire [(5'h11):(1'h0)] wire33;
  input wire signed [(4'h8):(1'h0)] wire32;
  input wire signed [(4'h8):(1'h0)] wire31;
  reg signed [(5'h10):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg66 = (1'h0);
  reg [(4'hf):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg62 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg61 = (1'h0);
  wire [(4'hd):(1'h0)] wire60;
  wire signed [(3'h6):(1'h0)] wire59;
  wire [(5'h13):(1'h0)] wire58;
  wire signed [(4'hc):(1'h0)] wire57;
  wire [(2'h2):(1'h0)] wire56;
  reg signed [(2'h2):(1'h0)] reg55 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg54 = (1'h0);
  reg [(5'h13):(1'h0)] reg53 = (1'h0);
  reg signed [(4'he):(1'h0)] reg52 = (1'h0);
  reg [(5'h11):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg50 = (1'h0);
  reg [(5'h13):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg47 = (1'h0);
  wire [(5'h15):(1'h0)] wire46;
  wire [(3'h4):(1'h0)] wire45;
  wire [(2'h2):(1'h0)] wire44;
  wire signed [(2'h3):(1'h0)] wire43;
  wire [(2'h3):(1'h0)] wire42;
  wire [(4'hc):(1'h0)] wire41;
  wire [(4'ha):(1'h0)] wire40;
  wire [(5'h12):(1'h0)] wire39;
  wire [(4'h9):(1'h0)] wire38;
  wire [(4'hd):(1'h0)] wire37;
  wire [(4'ha):(1'h0)] wire36;
  assign y = {reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 wire56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 wire42,
                 wire41,
                 wire40,
                 wire39,
                 wire38,
                 wire37,
                 wire36,
                 (1'h0)};
  assign wire36 = wire32;
  assign wire37 = wire32[(3'h7):(3'h6)];
  assign wire38 = (8'h9d);
  assign wire39 = wire32;
  assign wire40 = {$unsigned(wire37)};
  assign wire41 = (($unsigned(((wire36 ~^ wire32) + wire40)) >= (wire35 && ((!wire31) ~^ wire38))) ?
                      $signed($signed(($unsigned((8'hac)) <= wire31[(2'h3):(1'h1)]))) : $signed($signed($signed(wire31))));
  assign wire42 = ({$unsigned({{(8'haa), wire32},
                          (8'haa)})} || $unsigned((^wire32)));
  assign wire43 = wire40;
  assign wire44 = $unsigned(wire39);
  assign wire45 = $signed((~&(~|{$signed(wire35), $unsigned((8'had))})));
  assign wire46 = ({(+wire39)} ^~ (+(8'haa)));
  always
    @(posedge clk) begin
      reg47 <= ($unsigned(wire35[(3'h6):(2'h3)]) || $signed(wire45));
      reg48 <= ($unsigned(wire42) ?
          $unsigned(wire33) : ($unsigned((~&wire44[(1'h1):(1'h0)])) ?
              wire33[(5'h11):(1'h0)] : (($signed((8'hac)) - (wire34 << wire44)) << (wire43[(1'h1):(1'h1)] ?
                  (wire34 ? wire34 : (7'h43)) : $unsigned(reg47)))));
      if ($signed((($signed({wire42,
          reg47}) != (~&(-wire40))) < $signed(wire35[(4'hf):(2'h3)]))))
        begin
          reg49 <= (wire46[(2'h2):(1'h1)] >>> wire45);
          reg50 <= (((($unsigned(wire41) ?
              (wire32 <= wire41) : wire43) & $signed($signed(reg47))) << (8'h9e)) | (wire36[(3'h5):(1'h1)] >= ($unsigned((wire38 && wire37)) ~^ (^~{wire33}))));
          reg51 <= $signed((reg49[(4'hb):(4'ha)] ^~ {(|$signed(reg47)),
              wire34[(2'h2):(1'h1)]}));
          if ($unsigned(reg47[(2'h2):(1'h1)]))
            begin
              reg52 <= (8'h9e);
              reg53 <= $signed(($unsigned($unsigned((wire39 ?
                  (8'hb1) : wire32))) <= (~&{$signed(wire35)})));
            end
          else
            begin
              reg52 <= $signed((~$signed($unsigned((wire31 == wire46)))));
              reg53 <= $unsigned({$unsigned({$signed(wire31),
                      wire33[(4'ha):(2'h2)]})});
              reg54 <= wire32;
            end
        end
      else
        begin
          reg49 <= $signed(reg48);
          if ({$signed(wire35[(5'h11):(4'hb)])})
            begin
              reg50 <= ((reg51[(4'hd):(3'h5)] ?
                  (7'h40) : $unsigned((((7'h41) ~^ wire31) >> reg51))) | (wire43 ?
                  $signed(reg49) : (wire32[(3'h4):(2'h2)] * $signed((wire37 ?
                      (8'hbd) : (8'ha7))))));
              reg51 <= reg53;
              reg52 <= wire43[(1'h0):(1'h0)];
              reg53 <= (~^wire31);
              reg54 <= ((&((wire46 ?
                  (reg54 ?
                      reg48 : wire45) : reg50[(3'h5):(1'h1)]) != $unsigned(reg49[(1'h0):(1'h0)]))) != ((~wire37[(4'h9):(2'h2)]) ?
                  (reg47 ?
                      ((|wire33) > (+wire44)) : wire34[(1'h0):(1'h0)]) : ((&(^~wire37)) && ((^reg53) ?
                      {wire37} : ((8'hb6) << wire45)))));
            end
          else
            begin
              reg50 <= ($unsigned((8'h9d)) - $signed((!{((8'ha2) <= (8'hac)),
                  $unsigned(wire36)})));
              reg51 <= (8'hb6);
            end
        end
      reg55 <= $unsigned(($unsigned((((8'hb9) ?
          wire42 : (8'hbf)) >= reg53[(2'h3):(2'h2)])) | wire38[(4'h8):(2'h2)]));
    end
  assign wire56 = (wire39[(2'h2):(2'h2)] ^~ (+wire42));
  assign wire57 = reg50[(2'h3):(1'h1)];
  assign wire58 = {wire32, wire39[(2'h2):(2'h2)]};
  assign wire59 = {reg48[(4'h8):(3'h7)]};
  assign wire60 = $unsigned(($signed((wire46 ^~ $signed(reg51))) ?
                      $unsigned($signed(wire58[(5'h11):(1'h0)])) : wire40[(4'h8):(1'h0)]));
  always
    @(posedge clk) begin
      reg61 <= ($signed($unsigned($signed((wire36 >>> wire34)))) - wire46);
      reg62 <= (($unsigned($signed(wire38[(2'h3):(1'h1)])) ?
          ((8'hbb) - (wire41[(1'h0):(1'h0)] && wire58)) : (^$signed((reg51 < (8'ha7))))) != $unsigned(wire58[(3'h7):(3'h6)]));
      reg63 <= (wire37 >= $unsigned((wire40 ?
          reg55[(1'h0):(1'h0)] : wire35[(4'h9):(2'h3)])));
      reg64 <= $unsigned(reg50[(3'h5):(1'h0)]);
      reg65 <= (({reg53[(4'hb):(3'h4)]} ?
          $signed($signed((wire42 <= reg55))) : reg50) ^~ $signed(wire38[(1'h1):(1'h1)]));
    end
  always
    @(posedge clk) begin
      reg66 <= wire41[(4'h8):(2'h2)];
      reg67 <= ((&wire41[(3'h7):(2'h3)]) ? $signed(reg47) : (reg61 | (8'hb2)));
    end
endmodule