(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param199 = ((8'ha8) ? ({{(~(8'had))}, (((8'hbf) << (8'hb1)) ? ((8'hba) ^~ (7'h42)) : ((8'ha7) ? (7'h41) : (8'haf)))} ? (((+(8'hbb)) ? ((8'h9c) ~^ (8'hbc)) : (~&(8'hb2))) > (8'hba)) : ({((8'hac) ? (8'haf) : (8'ha4)), ((8'ha1) ? (8'hab) : (8'hbe))} ? (((8'hba) ? (8'hbc) : (7'h42)) ? ((8'ha4) ? (8'haa) : (8'ha1)) : ((8'ha0) ^~ (8'hb1))) : ({(8'ha5)} ? (^~(8'ha3)) : ((8'hba) == (8'ha1))))) : {((((8'hbb) - (8'hb6)) ^~ (~|(8'hbb))) ? (((8'haf) ? (8'ha0) : (8'ha6)) != ((7'h44) || (7'h40))) : (&((8'hb1) ? (8'h9c) : (8'hab)))), (-(!{(8'ha7), (8'hb7)}))})
, parameter param200 = (param199 >>> ((~&param199) && (8'h9e))) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1f4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire4;
  input wire signed [(4'h9):(1'h0)] wire3;
  input wire signed [(4'he):(1'h0)] wire2;
  input wire [(5'h10):(1'h0)] wire1;
  input wire [(5'h11):(1'h0)] wire0;
  wire [(4'hf):(1'h0)] wire198;
  reg signed [(4'h8):(1'h0)] reg197 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg196 = (1'h0);
  wire [(4'he):(1'h0)] wire195;
  wire [(3'h6):(1'h0)] wire194;
  reg [(4'hb):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg189 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg188 = (1'h0);
  reg [(3'h4):(1'h0)] reg187 = (1'h0);
  reg [(4'h8):(1'h0)] reg186 = (1'h0);
  reg [(4'ha):(1'h0)] reg185 = (1'h0);
  reg [(4'hc):(1'h0)] reg184 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg183 = (1'h0);
  reg [(5'h12):(1'h0)] reg182 = (1'h0);
  reg [(5'h13):(1'h0)] reg181 = (1'h0);
  reg [(2'h3):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg179 = (1'h0);
  reg [(4'hb):(1'h0)] reg178 = (1'h0);
  wire [(5'h10):(1'h0)] wire176;
  wire signed [(3'h5):(1'h0)] wire34;
  reg signed [(3'h6):(1'h0)] reg33 = (1'h0);
  reg [(3'h4):(1'h0)] reg32 = (1'h0);
  wire [(4'he):(1'h0)] wire31;
  wire signed [(4'h8):(1'h0)] wire30;
  wire signed [(4'hc):(1'h0)] wire29;
  wire signed [(4'ha):(1'h0)] wire28;
  reg signed [(3'h7):(1'h0)] reg27 = (1'h0);
  reg [(4'hf):(1'h0)] reg26 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg25 = (1'h0);
  reg [(4'hb):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg23 = (1'h0);
  reg [(5'h15):(1'h0)] reg22 = (1'h0);
  reg [(4'hc):(1'h0)] reg21 = (1'h0);
  reg [(4'h9):(1'h0)] reg20 = (1'h0);
  reg [(3'h4):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg18 = (1'h0);
  reg [(4'hd):(1'h0)] reg17 = (1'h0);
  reg signed [(4'he):(1'h0)] reg16 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg15 = (1'h0);
  reg [(4'hc):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg13 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg12 = (1'h0);
  reg [(2'h3):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg10 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire9;
  wire signed [(4'h8):(1'h0)] wire8;
  wire [(5'h12):(1'h0)] wire7;
  wire [(4'hc):(1'h0)] wire6;
  wire signed [(3'h4):(1'h0)] wire5;
  assign y = {wire198,
                 reg197,
                 reg196,
                 wire195,
                 wire194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 wire176,
                 wire34,
                 reg33,
                 reg32,
                 wire31,
                 wire30,
                 wire29,
                 wire28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 wire9,
                 wire8,
                 wire7,
                 wire6,
                 wire5,
                 (1'h0)};
  assign wire5 = $unsigned((+{((8'hb5) ? ((8'hab) < wire2) : $signed(wire2))}));
  assign wire6 = $signed(wire2);
  assign wire7 = wire6[(4'ha):(1'h0)];
  assign wire8 = (wire7[(3'h6):(2'h3)] ?
                     (+(~^wire2[(4'hd):(1'h1)])) : ($unsigned(wire0) < $signed($signed($unsigned(wire5)))));
  assign wire9 = (($unsigned(((^wire0) >>> $signed(wire6))) < wire6[(4'h9):(1'h1)]) != {($unsigned($signed(wire6)) ?
                         wire6[(4'hc):(3'h4)] : wire8)});
  always
    @(posedge clk) begin
      if ($signed($signed($signed($unsigned($signed(wire5))))))
        begin
          reg10 <= (|wire7);
          if (wire1[(4'hb):(2'h3)])
            begin
              reg11 <= wire2;
              reg12 <= wire0;
              reg13 <= $signed({($unsigned(wire2[(2'h3):(1'h0)]) + (~$unsigned(reg11)))});
            end
          else
            begin
              reg11 <= $unsigned(reg12[(3'h6):(3'h6)]);
              reg12 <= ({$unsigned($signed(wire1[(1'h0):(1'h0)]))} ?
                  (((^~wire9) & reg11) ?
                      $signed((|$signed(wire0))) : (($signed(wire6) && $signed(wire1)) - {(reg11 & (8'ha2)),
                          (-reg12)})) : ($signed(wire3[(2'h2):(2'h2)]) ?
                      wire7[(4'he):(4'hb)] : ((((8'ha1) ^~ wire4) | (~(8'hb4))) == $signed(reg12[(3'h7):(3'h4)]))));
              reg13 <= (8'hba);
              reg14 <= $signed($unsigned(($unsigned((reg13 == wire7)) ?
                  {(|(8'hb6)), $unsigned(reg11)} : (wire6[(4'ha):(4'h9)] ?
                      reg13[(2'h2):(1'h0)] : (!wire6)))));
              reg15 <= (^$unsigned($signed((8'had))));
            end
          reg16 <= reg14;
          reg17 <= $unsigned((-(^~$unsigned((wire3 ? (7'h42) : reg12)))));
          reg18 <= {wire8,
              $unsigned($unsigned(($unsigned(wire2) ?
                  $unsigned(wire8) : $unsigned(reg12))))};
        end
      else
        begin
          reg10 <= $signed({$unsigned((reg12[(3'h6):(1'h1)] ?
                  $signed((8'ha9)) : $signed(wire6)))});
          reg11 <= (~|($signed((~$signed(reg13))) ?
              $signed($signed($unsigned(reg18))) : reg18));
          reg12 <= $signed((^~reg13));
          reg13 <= ((!(~&reg12)) + (~|wire5[(1'h0):(1'h0)]));
        end
      reg19 <= ((~|{wire5[(2'h3):(2'h2)]}) != $unsigned(($unsigned((wire6 ?
              wire6 : wire7)) ?
          wire9 : $signed(wire9[(4'h9):(4'h9)]))));
      if ((!$unsigned(($signed(reg13) ?
          ((reg19 ? reg10 : (8'h9d)) ?
              wire3[(1'h1):(1'h0)] : reg11) : reg10[(1'h0):(1'h0)]))))
        begin
          reg20 <= $signed(wire8);
          reg21 <= (((wire7 * $signed(((8'hb9) << wire2))) ?
                  (^~$signed((reg18 ? wire9 : (8'had)))) : {(~^((8'hae) ?
                          wire3 : wire3))}) ?
              $signed(((~((8'hbb) ? reg17 : wire1)) ?
                  ({wire0} != (|reg18)) : wire4)) : $signed($signed((&(wire1 ?
                  wire9 : wire0)))));
          if ($signed($signed(($signed($unsigned((8'ha8))) || $signed({reg12})))))
            begin
              reg22 <= $signed(((&{(~^reg17), wire1}) ?
                  $signed($unsigned({reg14, reg14})) : $signed((-{reg14,
                      (8'ha4)}))));
            end
          else
            begin
              reg22 <= ($unsigned($signed(reg15)) ?
                  $signed(wire3) : $unsigned((~^$unsigned((wire8 ?
                      reg20 : reg14)))));
            end
        end
      else
        begin
          reg20 <= $signed(($signed((^~(!reg21))) ?
              (~&wire8[(2'h3):(2'h3)]) : $signed(wire0[(4'hc):(4'h9)])));
          if ($unsigned($unsigned(({(!reg15)} ?
              $unsigned($unsigned((8'haa))) : (~(reg17 ? (8'hb4) : wire2))))))
            begin
              reg21 <= {$unsigned($signed({(!wire5)}))};
              reg22 <= wire2;
              reg23 <= (reg15 ^~ $unsigned((|wire0[(4'h8):(3'h5)])));
              reg24 <= (!$signed(((&(wire4 ? reg16 : reg13)) ?
                  (((8'h9e) >= wire9) ?
                      (-(8'hbf)) : wire9[(1'h1):(1'h1)]) : $signed((|reg11)))));
              reg25 <= (reg21[(2'h3):(2'h2)] ?
                  (+(-((reg10 ?
                      wire2 : wire9) != (!(8'ha8))))) : {($unsigned((!reg12)) ?
                          {reg20} : ((reg11 ^ (8'hb4)) >>> ((8'ha8) | wire7))),
                      reg21[(2'h2):(1'h1)]});
            end
          else
            begin
              reg21 <= (+reg12);
              reg22 <= $unsigned($unsigned((($unsigned((8'hb5)) ?
                  (wire9 ? reg19 : wire6) : reg15) | wire4[(4'h8):(3'h5)])));
            end
          reg26 <= (($signed((+reg17[(3'h6):(1'h0)])) ?
              {($signed((8'hb0)) ?
                      reg24 : reg17)} : wire0) <= (!$unsigned((wire2 ?
              {wire3} : $signed(reg22)))));
          reg27 <= ((!$unsigned({$signed((8'hb5))})) ~^ ((~($signed(reg13) ?
              $unsigned(reg25) : $signed(reg26))) + reg19));
        end
    end
  assign wire28 = wire1[(4'hd):(1'h0)];
  assign wire29 = $signed((|reg18));
  assign wire30 = reg15;
  assign wire31 = reg19[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg32 <= ($signed((reg16[(3'h4):(1'h1)] && wire2[(4'ha):(1'h0)])) ?
          wire6 : $signed((8'hbf)));
      reg33 <= reg26;
    end
  assign wire34 = (~|$signed(reg15));
  module35 modinst177 (wire176, clk, wire0, wire31, wire1, wire7);
  always
    @(posedge clk) begin
      reg178 <= (~|(wire8 >> reg27[(2'h3):(2'h2)]));
      reg179 <= (wire5 ?
          reg13 : (({(!wire176)} ?
              (((8'hac) <<< wire7) ?
                  wire29 : (reg22 ?
                      reg13 : reg12)) : reg23[(2'h2):(1'h1)]) + $unsigned(reg32)));
      if (({reg26, (~({wire9} ? (wire7 <<< reg13) : reg24[(1'h1):(1'h0)]))} ?
          (($unsigned(reg19[(2'h2):(1'h0)]) <= wire176[(4'he):(4'h8)]) ?
              $unsigned($unsigned(reg10[(1'h0):(1'h0)])) : (!($unsigned(wire2) << (reg179 <= wire34)))) : reg14[(2'h2):(1'h0)]))
        begin
          reg180 <= $signed(reg11);
          if (wire9)
            begin
              reg181 <= $unsigned(($signed({$signed(reg25),
                      (wire34 ? reg178 : (8'ha7))}) ?
                  ((^~$unsigned(reg24)) ?
                      $signed((+reg21)) : wire0) : reg17[(4'ha):(3'h7)]));
              reg182 <= (~|((~&wire5[(1'h1):(1'h0)]) >= reg13));
              reg183 <= (reg10[(3'h5):(3'h5)] | wire31);
              reg184 <= (reg14[(3'h5):(2'h3)] ?
                  (8'h9f) : (reg11[(2'h2):(2'h2)] <= {$signed(reg10),
                      (+(8'hab))}));
            end
          else
            begin
              reg181 <= $signed($signed({$unsigned({reg27, reg178}),
                  $unsigned(wire9)}));
              reg182 <= (reg14 ?
                  $signed(reg181) : $unsigned((reg23[(3'h4):(2'h3)] ?
                      $signed($signed(reg23)) : reg27[(1'h1):(1'h0)])));
            end
          reg185 <= (^wire34[(3'h5):(3'h5)]);
        end
      else
        begin
          reg180 <= $unsigned((wire8[(1'h1):(1'h0)] << wire2[(4'h9):(3'h6)]));
          reg181 <= (~^wire28);
          reg182 <= ($unsigned((~&reg180[(1'h1):(1'h0)])) >> $signed({reg13[(2'h3):(2'h2)],
              wire4[(4'hb):(3'h7)]}));
        end
      if (($unsigned(reg20[(3'h7):(3'h5)]) ~^ $signed(($signed($signed(reg32)) <<< reg23))))
        begin
          reg186 <= $unsigned(({$unsigned(reg183[(1'h1):(1'h1)]),
                  $signed((wire31 << reg25))} ?
              reg23 : ((((8'ha5) ? reg10 : reg22) ?
                  $signed(reg15) : $unsigned(wire31)) != {(wire9 + reg11)})));
          reg187 <= $signed((reg16 & $signed((reg26 >> (reg25 <<< reg178)))));
          reg188 <= reg27;
          if (($signed(($signed((wire28 * reg13)) ?
                  $unsigned($signed(reg27)) : $signed({(8'ha3)}))) ?
              (^$unsigned({(reg22 ? wire31 : reg182),
                  $signed(reg17)})) : (&(reg16[(4'hb):(4'ha)] ?
                  $unsigned($unsigned(reg180)) : (~^(!reg13))))))
            begin
              reg189 <= $signed((reg183 >> ({reg18} < ((reg179 - reg17) ?
                  reg12[(1'h1):(1'h0)] : $signed(wire2)))));
              reg190 <= {($signed(reg14[(2'h2):(1'h1)]) <<< reg24)};
              reg191 <= $unsigned((($signed({reg178, (7'h43)}) ?
                      reg181 : (+(reg16 ? reg32 : (8'hbf)))) ?
                  reg178[(1'h0):(1'h0)] : $unsigned($signed((reg17 > wire34)))));
            end
          else
            begin
              reg189 <= (-$signed((+reg188)));
              reg190 <= $signed($signed(reg15));
              reg191 <= reg14[(4'h9):(4'h9)];
              reg192 <= $signed((((wire28 ? reg14[(1'h1):(1'h0)] : (^reg179)) ?
                      $signed($unsigned(reg33)) : $unsigned((reg20 ?
                          (8'hb9) : (8'h9c)))) ?
                  (|(reg32[(1'h0):(1'h0)] ?
                      (reg11 < reg179) : $signed(wire8))) : ($unsigned($signed(wire6)) << reg183[(2'h2):(1'h0)])));
              reg193 <= (((($unsigned(reg15) <<< $unsigned(reg190)) <= (wire6[(3'h7):(2'h3)] >>> (reg13 == reg12))) != reg185[(4'ha):(4'h8)]) * ($unsigned($unsigned(wire176[(4'hb):(1'h0)])) | $signed(reg23[(2'h2):(2'h2)])));
            end
        end
      else
        begin
          reg186 <= (wire4[(4'hf):(4'hc)] ?
              (~|{$signed((8'hac))}) : ((|((&reg180) | (-reg179))) ?
                  reg186 : ((wire6 < (~&reg23)) == reg192)));
        end
    end
  assign wire194 = wire3[(1'h1):(1'h0)];
  assign wire195 = $signed((-$unsigned(reg32[(1'h1):(1'h1)])));
  always
    @(posedge clk) begin
      reg196 <= ($unsigned((($signed(reg191) || $unsigned(wire194)) & (reg183[(2'h2):(1'h0)] ?
          $signed(reg191) : (reg189 ?
              wire30 : reg26)))) >> reg189[(3'h4):(3'h4)]);
      reg197 <= (8'hbe);
    end
  assign wire198 = (!(+(($unsigned(wire9) ?
                       $signed(reg14) : $signed(reg193)) == {(^(8'hb7)),
                       (wire195 ? wire1 : (8'h9d))})));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module35
#( parameter param174 = ((((~&(!(7'h42))) <<< (((8'hbc) ? (8'hb2) : (8'ha4)) ? {(8'hb0), (8'ha6)} : {(8'hbf)})) ? ({{(8'ha0)}} ~^ ((!(7'h44)) ? ((8'hb9) ? (8'hb7) : (8'ha8)) : ((7'h40) ? (8'ha8) : (8'hb6)))) : ((((8'ha6) ^ (8'hb2)) | ((8'hb8) != (8'ha6))) <<< ((|(8'ha5)) ? ((8'hb5) ? (7'h44) : (8'had)) : {(8'h9f), (8'ha0)}))) < (((((8'ha1) ^~ (8'ha5)) ? (~^(8'ha8)) : {(8'hbc)}) | (((8'h9e) ? (8'hb2) : (8'hbd)) + {(8'h9d)})) ^ ((((8'hb4) && (7'h41)) >>> ((8'hb4) ? (7'h41) : (8'ha0))) || (((7'h44) > (8'h9f)) ? ((8'hbe) ? (8'h9e) : (8'hbf)) : {(8'hb7)}))))
, parameter param175 = {{({(-param174)} <= (param174 | (param174 & param174))), (8'hb3)}} )
(y, clk, wire36, wire37, wire38, wire39);
  output wire [(32'h12d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire36;
  input wire [(4'he):(1'h0)] wire37;
  input wire [(4'hc):(1'h0)] wire38;
  input wire [(4'hf):(1'h0)] wire39;
  wire signed [(5'h15):(1'h0)] wire173;
  wire [(5'h14):(1'h0)] wire172;
  wire signed [(4'he):(1'h0)] wire170;
  wire [(2'h3):(1'h0)] wire155;
  wire [(5'h10):(1'h0)] wire154;
  reg signed [(5'h15):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg42 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg43 = (1'h0);
  reg [(5'h12):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg45 = (1'h0);
  reg [(3'h7):(1'h0)] reg46 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg47 = (1'h0);
  reg [(5'h12):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg49 = (1'h0);
  reg [(5'h13):(1'h0)] reg50 = (1'h0);
  reg [(3'h5):(1'h0)] reg51 = (1'h0);
  reg [(5'h11):(1'h0)] reg52 = (1'h0);
  reg signed [(4'he):(1'h0)] reg53 = (1'h0);
  reg [(4'hc):(1'h0)] reg54 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg55 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire83;
  wire signed [(3'h7):(1'h0)] wire152;
  assign y = {wire173,
                 wire172,
                 wire170,
                 wire155,
                 wire154,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 reg54,
                 reg55,
                 wire83,
                 wire152,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((($signed(wire38) || $unsigned(wire36)) ?
          {$unsigned((wire37 >>> (wire38 ?
                  wire39 : wire36)))} : $signed({((|wire36) ?
                  (wire36 ? wire36 : wire39) : wire39),
              (^{wire38})})))
        begin
          reg40 <= (+wire39);
          reg41 <= ($signed($signed($unsigned((!wire37)))) ?
              $signed(reg40[(5'h15):(2'h3)]) : wire36[(4'h8):(3'h5)]);
        end
      else
        begin
          reg40 <= $signed((^wire39[(4'h9):(2'h3)]));
          if ($unsigned(wire36))
            begin
              reg41 <= $unsigned(((+reg40[(4'hb):(1'h1)]) || $signed((|$unsigned(wire39)))));
              reg42 <= ((8'hbd) == $signed($signed(wire38[(3'h5):(1'h0)])));
              reg43 <= (reg42[(5'h10):(4'he)] <<< $unsigned((wire38 ?
                  {(wire39 ? reg40 : (8'haf)), $unsigned(wire37)} : (8'ha4))));
              reg44 <= $signed((!(~$signed({reg43, reg40}))));
              reg45 <= ((+$unsigned(wire39)) >> $unsigned(({$unsigned(reg40),
                      wire36} ?
                  ($unsigned(wire36) ^ (8'haf)) : ($signed(wire39) ?
                      reg41 : (-wire36)))));
            end
          else
            begin
              reg41 <= reg40[(3'h4):(1'h0)];
              reg42 <= (~^$signed((((wire37 < wire36) && (~|reg40)) ?
                  reg44[(3'h5):(1'h1)] : ((wire38 ?
                      wire37 : wire39) - (^~reg40)))));
            end
          if (wire37)
            begin
              reg46 <= reg45;
              reg47 <= reg45;
            end
          else
            begin
              reg46 <= ((~^$unsigned((~|(!reg44)))) && (((-$unsigned(wire38)) >>> wire37) ?
                  wire36[(2'h2):(1'h1)] : (wire37 >> $unsigned((reg47 == reg43)))));
              reg47 <= (8'haf);
              reg48 <= $unsigned(reg46[(2'h3):(2'h3)]);
              reg49 <= (7'h43);
              reg50 <= reg41[(2'h3):(2'h2)];
            end
        end
      if (((wire37[(2'h2):(2'h2)] > wire38) ?
          reg40 : (reg42 ?
              ({$signed(reg40), (reg40 == reg40)} >>> (wire38[(3'h4):(3'h4)] ?
                  (+(8'hac)) : wire37)) : reg49[(4'hc):(3'h4)])))
        begin
          reg51 <= ($signed(((|(wire37 && reg45)) ?
              {reg42[(5'h13):(4'he)]} : $signed((reg49 ?
                  reg45 : reg44)))) * $signed($unsigned($unsigned($signed(wire39)))));
          reg52 <= ((8'had) ?
              (&reg46[(2'h2):(2'h2)]) : $signed(($signed($signed(wire36)) >> {(reg45 >> reg49)})));
          reg53 <= ((wire37 < reg51[(2'h2):(2'h2)]) ?
              $signed($unsigned(reg41[(3'h5):(1'h1)])) : wire37);
        end
      else
        begin
          reg51 <= reg52[(2'h2):(1'h0)];
          reg52 <= {$unsigned($signed($signed({reg40})))};
          reg53 <= $signed((~&$unsigned($signed($unsigned(reg49)))));
          reg54 <= (((($unsigned(reg53) ?
              $unsigned(reg46) : (&wire38)) == reg47[(3'h6):(1'h0)]) & ((reg42[(5'h10):(3'h6)] ?
                  $unsigned(reg49) : (-reg53)) ?
              ($signed(reg48) ?
                  reg43 : reg47) : (~&reg42[(3'h7):(3'h4)]))) ^ (-$signed(((reg48 ^~ wire39) >>> $signed(reg52)))));
        end
      reg55 <= reg46[(1'h1):(1'h0)];
    end
  module56 modinst84 (.wire58(reg42), .wire59(wire37), .clk(clk), .wire57(reg55), .y(wire83), .wire60(reg41));
  module85 modinst153 (.wire89(reg45), .y(wire152), .wire90(wire39), .wire86(reg41), .clk(clk), .wire87(reg44), .wire88(reg47));
  assign wire154 = (!{$signed(((~&wire36) <<< {reg53, wire83})),
                       (reg45[(3'h6):(3'h6)] << (-{wire38}))});
  assign wire155 = (8'hbb);
  module156 modinst171 (wire170, clk, wire38, reg50, reg43, wire83);
  assign wire172 = $signed({reg55,
                       $signed({$signed(reg55), (reg50 ? (8'had) : wire170)})});
  assign wire173 = wire37[(4'hc):(4'hc)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module156  (y, clk, wire160, wire159, wire158, wire157);
  output wire [(32'h5a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire160;
  input wire [(4'hb):(1'h0)] wire159;
  input wire signed [(2'h2):(1'h0)] wire158;
  input wire [(4'h8):(1'h0)] wire157;
  wire signed [(4'hc):(1'h0)] wire169;
  wire signed [(2'h2):(1'h0)] wire168;
  reg [(3'h7):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg166 = (1'h0);
  wire [(5'h10):(1'h0)] wire165;
  wire [(3'h6):(1'h0)] wire164;
  wire signed [(3'h7):(1'h0)] wire163;
  wire signed [(4'hc):(1'h0)] wire162;
  wire [(4'hb):(1'h0)] wire161;
  assign y = {wire169,
                 wire168,
                 reg167,
                 reg166,
                 wire165,
                 wire164,
                 wire163,
                 wire162,
                 wire161,
                 (1'h0)};
  assign wire161 = (8'hbf);
  assign wire162 = ($signed(wire157[(2'h3):(2'h2)]) ~^ $unsigned({wire160[(4'ha):(1'h1)],
                       {wire161[(2'h2):(2'h2)]}}));
  assign wire163 = ($signed($signed(((wire161 ^ wire162) || $signed((8'hb5))))) ?
                       $signed((wire160 ?
                           ({wire159, wire157} | (wire162 ?
                               wire157 : wire157)) : ((wire159 >= wire160) ?
                               $unsigned(wire157) : wire160[(1'h1):(1'h0)]))) : wire159);
  assign wire164 = {(wire157 ~^ wire157[(3'h6):(2'h2)]), (!wire160)};
  assign wire165 = (-$unsigned(wire162[(4'ha):(3'h5)]));
  always
    @(posedge clk) begin
      reg166 <= wire163[(1'h1):(1'h0)];
      reg167 <= wire157;
    end
  assign wire168 = {reg166};
  assign wire169 = $unsigned(wire157[(3'h4):(2'h2)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module85
#( parameter param151 = {(~|((~{(8'ha8)}) != (^((8'ha9) ? (8'ha3) : (8'h9f))))), (7'h40)} )
(y, clk, wire90, wire89, wire88, wire87, wire86);
  output wire [(32'h2ab):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire90;
  input wire signed [(3'h7):(1'h0)] wire89;
  input wire [(4'h8):(1'h0)] wire88;
  input wire signed [(5'h12):(1'h0)] wire87;
  input wire [(2'h2):(1'h0)] wire86;
  wire signed [(4'hd):(1'h0)] wire150;
  wire signed [(3'h7):(1'h0)] wire149;
  wire [(3'h5):(1'h0)] wire148;
  wire [(3'h6):(1'h0)] wire147;
  reg [(2'h2):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg145 = (1'h0);
  wire [(5'h13):(1'h0)] wire144;
  wire [(3'h5):(1'h0)] wire143;
  wire signed [(5'h10):(1'h0)] wire142;
  wire [(5'h10):(1'h0)] wire141;
  wire [(2'h3):(1'h0)] wire140;
  wire [(4'he):(1'h0)] wire139;
  wire signed [(5'h10):(1'h0)] wire138;
  reg [(3'h4):(1'h0)] reg137 = (1'h0);
  reg signed [(4'he):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg132 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg129 = (1'h0);
  reg [(4'h8):(1'h0)] reg128 = (1'h0);
  reg [(4'he):(1'h0)] reg127 = (1'h0);
  reg [(3'h6):(1'h0)] reg126 = (1'h0);
  reg [(5'h12):(1'h0)] reg125 = (1'h0);
  reg [(4'hf):(1'h0)] reg124 = (1'h0);
  reg [(4'hc):(1'h0)] reg123 = (1'h0);
  reg [(4'h9):(1'h0)] reg122 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg121 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg120 = (1'h0);
  reg [(4'hf):(1'h0)] reg119 = (1'h0);
  reg [(4'ha):(1'h0)] reg118 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire117;
  wire signed [(4'h8):(1'h0)] wire116;
  wire [(4'hd):(1'h0)] wire115;
  reg [(3'h6):(1'h0)] reg114 = (1'h0);
  reg [(4'he):(1'h0)] reg113 = (1'h0);
  reg [(4'h8):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg111 = (1'h0);
  reg [(4'h9):(1'h0)] reg110 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire109;
  wire [(5'h12):(1'h0)] wire108;
  wire signed [(5'h12):(1'h0)] wire107;
  reg [(3'h4):(1'h0)] reg106 = (1'h0);
  reg [(4'hc):(1'h0)] reg105 = (1'h0);
  reg [(4'hf):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg103 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg101 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg100 = (1'h0);
  reg [(5'h12):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg98 = (1'h0);
  reg [(4'hb):(1'h0)] reg97 = (1'h0);
  reg [(4'he):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg95 = (1'h0);
  reg [(4'he):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg93 = (1'h0);
  wire [(3'h7):(1'h0)] wire92;
  wire signed [(4'h9):(1'h0)] wire91;
  assign y = {wire150,
                 wire149,
                 wire148,
                 wire147,
                 reg146,
                 reg145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 wire117,
                 wire116,
                 wire115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 wire109,
                 wire108,
                 wire107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 wire92,
                 wire91,
                 (1'h0)};
  assign wire91 = wire86;
  assign wire92 = wire86[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      if (wire91)
        begin
          reg93 <= (((+$unsigned($signed(wire88))) | {wire87[(4'he):(4'he)],
                  (wire89[(3'h4):(2'h2)] ? $signed(wire86) : wire86)}) ?
              wire87[(4'ha):(3'h4)] : $unsigned(wire88));
          if (wire91)
            begin
              reg94 <= $unsigned((~|(wire86[(1'h0):(1'h0)] ?
                  reg93[(1'h1):(1'h1)] : {{wire88}})));
              reg95 <= wire86;
              reg96 <= wire92[(1'h1):(1'h0)];
            end
          else
            begin
              reg94 <= reg94[(3'h6):(3'h5)];
              reg95 <= wire92[(3'h4):(3'h4)];
              reg96 <= reg93;
              reg97 <= (8'hbd);
            end
          reg98 <= {(-reg93)};
        end
      else
        begin
          reg93 <= wire86;
          reg94 <= wire92[(3'h7):(3'h6)];
          reg95 <= $signed({(reg98 >>> (-(reg96 ? reg98 : reg98))),
              $signed(($unsigned(wire91) ?
                  $unsigned(reg94) : $unsigned(reg96)))});
          reg96 <= wire87;
          reg97 <= (-wire88[(3'h4):(2'h3)]);
        end
      if (($signed(((-$signed(wire92)) <= ((reg94 ? (8'hb1) : reg98) ?
          (reg97 >= wire92) : $unsigned(wire87)))) <<< reg95))
        begin
          reg99 <= wire86[(2'h2):(1'h1)];
          reg100 <= reg98;
          if (((+$unsigned(((^~wire92) > wire87))) - $unsigned($unsigned(wire90[(3'h6):(3'h5)]))))
            begin
              reg101 <= (reg98 ?
                  wire87[(4'h9):(1'h1)] : ((-(^wire90)) == (&wire92)));
              reg102 <= $unsigned($signed(((~|reg100[(1'h1):(1'h0)]) ?
                  ((~|wire87) ~^ wire92) : ($signed(wire86) << (reg97 ?
                      reg101 : wire91)))));
            end
          else
            begin
              reg101 <= reg94;
              reg102 <= (&(|(|($unsigned((8'hb0)) ?
                  ((8'hbc) ? reg98 : wire87) : reg93[(4'hc):(4'hc)]))));
              reg103 <= (|wire89[(3'h5):(3'h5)]);
              reg104 <= $unsigned((wire91 ?
                  ($unsigned((reg93 & (8'hb4))) * reg94[(2'h3):(2'h3)]) : reg95));
              reg105 <= ($signed((&wire87[(1'h0):(1'h0)])) < ((reg101 ?
                  wire91[(1'h0):(1'h0)] : ((^~reg100) >>> (~|wire89))) ^~ (^~reg96[(4'he):(3'h4)])));
            end
        end
      else
        begin
          reg99 <= (8'h9d);
        end
      if (((~$signed($unsigned((reg103 ?
          reg101 : wire86)))) || (reg93 << reg99[(1'h0):(1'h0)])))
        begin
          reg106 <= $signed((~&(^~{$signed(reg94)})));
        end
      else
        begin
          reg106 <= ($unsigned({(~(^~wire88)),
              ((wire89 ?
                  reg102 : reg96) ~^ $unsigned(reg104))}) ^~ wire87[(1'h0):(1'h0)]);
        end
    end
  assign wire107 = $signed($signed((wire88 ?
                       $signed(wire90[(1'h0):(1'h0)]) : $unsigned({(8'hb6),
                           (8'h9d)}))));
  assign wire108 = $signed((reg93[(4'hc):(4'ha)] ?
                       ((8'hb8) ?
                           (|{reg99}) : (wire107[(5'h10):(4'he)] ~^ wire107)) : reg96[(2'h3):(2'h3)]));
  assign wire109 = {reg100};
  always
    @(posedge clk) begin
      reg110 <= reg104[(3'h7):(1'h0)];
      reg111 <= $signed(((~(wire89[(3'h5):(2'h2)] ? reg105 : wire87)) ?
          ((~(~^reg99)) ?
              $signed($unsigned((8'hbc))) : (~^{wire90})) : reg105));
      if ({$unsigned((($signed(wire107) <= (reg97 * wire86)) < (^$signed((8'hb5))))),
          $unsigned(((&(wire109 ~^ wire88)) ?
              ($signed(reg95) + $unsigned(reg95)) : $signed(reg104)))})
        begin
          reg112 <= (~$unsigned(reg111[(1'h1):(1'h0)]));
          reg113 <= (+{wire86[(2'h2):(1'h1)]});
        end
      else
        begin
          reg112 <= (reg111 ?
              reg100 : ($signed($unsigned((reg98 <= reg110))) ?
                  (((+wire87) ? (reg95 >>> reg110) : (-reg104)) ?
                      (!(|(8'h9d))) : wire107[(2'h3):(2'h2)]) : reg96[(4'he):(3'h6)]));
          reg113 <= reg100[(1'h1):(1'h0)];
          reg114 <= $signed(reg95[(2'h3):(2'h2)]);
        end
    end
  assign wire115 = ((wire108 ?
                           {$signed({wire89}),
                               ($unsigned(reg102) ?
                                   (reg114 ?
                                       wire108 : reg97) : {reg102})} : {reg103}) ?
                       (-$unsigned({{wire109, wire89},
                           reg100[(2'h2):(1'h1)]})) : reg105[(4'hb):(4'hb)]);
  assign wire116 = $signed(($unsigned(wire108) ?
                       ({(reg114 ? reg110 : reg111),
                               (reg111 ? wire89 : reg97)} ?
                           (reg105[(3'h5):(2'h3)] ?
                               $signed(reg97) : $unsigned((8'hba))) : (-wire109)) : (+$unsigned(reg100[(1'h1):(1'h0)]))));
  assign wire117 = ($unsigned(((reg100[(1'h1):(1'h0)] ?
                           wire115 : reg93[(3'h5):(2'h2)]) != {reg96,
                           $signed(reg103)})) ?
                       (wire108[(3'h6):(3'h6)] ?
                           reg103[(3'h4):(1'h1)] : {{(8'hb4),
                                   (~reg113)}}) : reg114);
  always
    @(posedge clk) begin
      reg118 <= ((wire86[(2'h2):(1'h0)] + $unsigned($unsigned($unsigned(reg99)))) <= reg95);
      reg119 <= ((|wire107) ?
          (!(&(+(wire116 ? reg103 : wire117)))) : (|(~(~{wire86, reg113}))));
      if ((+$unsigned(($unsigned(reg97[(3'h6):(3'h5)]) ?
          $signed(reg98[(4'he):(4'ha)]) : ((reg99 ?
              reg94 : wire117) >>> (wire115 + reg103))))))
        begin
          reg120 <= $signed(reg112[(3'h4):(2'h2)]);
          reg121 <= (reg101 ?
              $signed((((~^reg97) ?
                  $signed(wire89) : ((8'ha8) >> (8'hb9))) < $signed(wire87[(4'ha):(3'h5)]))) : reg93[(1'h1):(1'h1)]);
          reg122 <= reg96[(3'h4):(3'h4)];
        end
      else
        begin
          if (((^~($signed((reg121 >> wire107)) < ($unsigned(reg113) ?
                  (wire108 ? reg105 : reg121) : (-wire109)))) ?
              {(^~$signed($signed(reg110)))} : reg96[(4'h8):(3'h6)]))
            begin
              reg120 <= (~^reg104);
              reg121 <= (~^(($unsigned(reg118) << {(wire115 ? reg114 : (8'h9d)),
                  reg111[(1'h1):(1'h1)]}) && (-$unsigned((!reg98)))));
            end
          else
            begin
              reg120 <= wire86[(1'h1):(1'h0)];
              reg121 <= reg103[(4'hc):(1'h0)];
              reg122 <= reg101;
            end
          reg123 <= (8'h9c);
          reg124 <= (+reg122[(2'h2):(1'h1)]);
          reg125 <= ((~$signed((~&wire90[(1'h1):(1'h1)]))) ?
              {$unsigned(reg119[(1'h1):(1'h1)])} : reg114);
          reg126 <= (8'ha9);
        end
      reg127 <= (((reg106 ? $unsigned(reg93) : (^~$unsigned(wire86))) ?
              reg102[(1'h0):(1'h0)] : {((reg126 ? reg99 : reg100) > (-wire109)),
                  $unsigned((~|reg94))}) ?
          wire116[(3'h4):(2'h2)] : $unsigned((((^wire108) ?
                  $unsigned(reg113) : (wire109 ? (8'hb1) : wire86)) ?
              reg101 : reg122)));
      if ({(reg97[(1'h0):(1'h0)] ? $signed(reg104[(4'hb):(3'h4)]) : (^reg104)),
          ((reg96 >>> ({(8'ha3), (8'hbe)} != reg96)) << wire92[(3'h5):(3'h5)])})
        begin
          reg128 <= reg120[(3'h4):(3'h4)];
          if ($unsigned($unsigned($unsigned($unsigned(wire116[(3'h4):(2'h3)])))))
            begin
              reg129 <= $unsigned(wire115);
            end
          else
            begin
              reg129 <= reg100[(2'h2):(1'h1)];
              reg130 <= reg124;
              reg131 <= $unsigned($signed((($signed((8'hbe)) >> $signed(wire87)) ?
                  $signed((8'hb0)) : wire108[(4'h8):(1'h1)])));
              reg132 <= reg128[(1'h1):(1'h1)];
            end
          if ($signed((-((~|reg125) ^~ (reg98[(4'hf):(3'h5)] ?
              (~&reg125) : $signed(reg100))))))
            begin
              reg133 <= reg124[(3'h5):(2'h2)];
              reg134 <= $signed(wire115);
              reg135 <= $signed(((($unsigned(wire86) ?
                      reg104 : (reg101 ? reg97 : reg121)) ?
                  $signed((&reg110)) : ((reg114 || wire115) ?
                      {wire115} : (&reg101))) > {$signed((reg121 ^ wire117)),
                  $signed((wire92 ? wire117 : reg99))}));
            end
          else
            begin
              reg133 <= reg105;
              reg134 <= (8'hbf);
              reg135 <= ($signed((!{$unsigned(wire86),
                  (reg121 + reg121)})) >> reg126);
            end
        end
      else
        begin
          if ({((+(~^$unsigned(wire107))) == wire86),
              {$signed((~^reg130[(4'h8):(1'h1)])), {(8'hae), {(^reg123)}}}})
            begin
              reg128 <= ((!$signed(({reg121} ?
                      ((8'ha9) ? (7'h42) : reg106) : {(8'ha2)}))) ?
                  $unsigned({reg135[(4'hb):(3'h5)]}) : $signed(reg119[(1'h0):(1'h0)]));
              reg129 <= reg113;
            end
          else
            begin
              reg128 <= $signed((!(wire92[(1'h0):(1'h0)] ?
                  reg105 : (reg99[(2'h3):(1'h0)] + wire92[(3'h7):(2'h3)]))));
              reg129 <= reg93[(5'h10):(3'h5)];
            end
          reg130 <= (-$unsigned($unsigned((8'haa))));
          reg131 <= $unsigned($unsigned(wire107));
          if ($signed($unsigned((-(^~{wire86})))))
            begin
              reg132 <= reg113;
              reg133 <= (((^~reg134[(2'h3):(2'h3)]) ?
                      (reg97[(1'h0):(1'h0)] < $signed($unsigned(reg127))) : (((~^reg123) >> $signed(reg104)) || reg105)) ?
                  (!(8'h9c)) : (reg95 ? wire107 : (reg98 < (-(8'hae)))));
              reg134 <= {wire115};
              reg135 <= ($unsigned(reg93[(4'hd):(3'h4)]) & reg118);
              reg136 <= ((^~reg103[(4'hc):(3'h4)]) >>> reg122);
            end
          else
            begin
              reg132 <= wire117;
            end
          reg137 <= ($signed((reg132 + $unsigned((reg124 <<< reg112)))) ?
              reg127 : ($signed({reg121}) ?
                  ($unsigned($unsigned(reg114)) + $signed($unsigned(reg113))) : (((&(8'hb4)) ?
                      (reg100 ? reg98 : reg103) : (reg130 ?
                          reg129 : (8'hb7))) >> (+((8'ha2) ?
                      reg111 : reg135)))));
        end
    end
  assign wire138 = ($unsigned($signed((8'hb2))) ?
                       reg137 : $unsigned((reg96[(2'h3):(1'h1)] == (~$unsigned(reg127)))));
  assign wire139 = $signed(((~|reg134) || $signed($signed($signed(wire115)))));
  assign wire140 = (!reg112[(3'h5):(1'h0)]);
  assign wire141 = ($signed(wire91[(4'h8):(3'h7)]) ?
                       (reg136 ?
                           reg103 : $unsigned(($signed(reg113) - reg121[(1'h0):(1'h0)]))) : {$unsigned($signed($unsigned((8'ha3))))});
  assign wire142 = {((reg98 != $unsigned($unsigned(reg112))) ?
                           ((+wire108) ?
                               {(reg104 > reg95)} : ($signed(wire139) == $unsigned(reg101))) : wire108),
                       (-(8'ha2))};
  assign wire143 = (reg122 ?
                       (((reg112 & (wire140 ? reg97 : (8'hac))) ?
                               ((~&(8'ha3)) ?
                                   (wire108 && reg129) : $unsigned((8'hbb))) : (^(~reg103))) ?
                           (!$unsigned($signed(reg97))) : (^($unsigned((8'ha6)) <<< (reg119 ?
                               (8'ha5) : reg123)))) : {((wire92[(3'h7):(3'h4)] ?
                                   (8'hb4) : (8'ha0)) ?
                               reg122[(3'h7):(1'h1)] : $signed((~^reg94)))});
  assign wire144 = (8'hb8);
  always
    @(posedge clk) begin
      reg145 <= ((8'hb4) > ((+$unsigned($unsigned((8'hbf)))) <= (~|$unsigned((reg113 + wire92)))));
      reg146 <= reg99[(3'h5):(3'h5)];
    end
  assign wire147 = reg119[(4'h9):(1'h1)];
  assign wire148 = (!$signed($unsigned((~^reg133[(3'h4):(2'h2)]))));
  assign wire149 = (($signed(reg101[(4'ha):(2'h3)]) ?
                           ($unsigned((wire108 || reg104)) >>> $unsigned(reg146[(1'h1):(1'h1)])) : reg97[(3'h7):(3'h6)]) ?
                       $unsigned(reg134[(1'h1):(1'h0)]) : $signed(reg103));
  assign wire150 = {($unsigned($unsigned($unsigned(reg125))) * $unsigned($signed({reg129})))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module56  (y, clk, wire60, wire59, wire58, wire57);
  output wire [(32'h11f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire60;
  input wire [(4'he):(1'h0)] wire59;
  input wire [(5'h14):(1'h0)] wire58;
  input wire [(2'h3):(1'h0)] wire57;
  wire [(4'hc):(1'h0)] wire82;
  wire signed [(4'hd):(1'h0)] wire81;
  wire [(4'hb):(1'h0)] wire80;
  wire signed [(3'h4):(1'h0)] wire79;
  wire signed [(5'h10):(1'h0)] wire78;
  wire [(4'h8):(1'h0)] wire77;
  wire [(4'hd):(1'h0)] wire76;
  wire [(4'hd):(1'h0)] wire75;
  wire [(4'h8):(1'h0)] wire74;
  wire [(3'h7):(1'h0)] wire73;
  wire signed [(5'h11):(1'h0)] wire72;
  wire [(4'ha):(1'h0)] wire71;
  wire signed [(4'ha):(1'h0)] wire70;
  wire [(5'h10):(1'h0)] wire69;
  wire signed [(5'h14):(1'h0)] wire68;
  wire [(4'h9):(1'h0)] wire67;
  wire signed [(4'hc):(1'h0)] wire66;
  wire [(5'h13):(1'h0)] wire65;
  wire signed [(5'h14):(1'h0)] wire64;
  wire [(4'hd):(1'h0)] wire63;
  wire signed [(5'h15):(1'h0)] wire62;
  wire [(4'he):(1'h0)] wire61;
  assign y = {wire82,
                 wire81,
                 wire80,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire74,
                 wire73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 (1'h0)};
  assign wire61 = (~&wire58);
  assign wire62 = $unsigned($unsigned((|$signed($unsigned(wire61)))));
  assign wire63 = wire61[(1'h0):(1'h0)];
  assign wire64 = (({wire57[(1'h1):(1'h0)]} ?
                          (({(8'ha6)} && $signed((8'had))) ?
                              ($signed((8'hbe)) ?
                                  wire57[(2'h3):(2'h3)] : (wire63 ^~ (7'h41))) : ($unsigned(wire62) ?
                                  (wire63 && wire57) : (wire61 <<< wire59))) : ((8'hb6) ?
                              wire57 : wire59[(4'he):(4'hb)])) ?
                      (~|wire58) : wire58);
  assign wire65 = $unsigned(((!$signed(wire59[(4'hd):(4'hb)])) ?
                      (&$signed((wire63 - wire63))) : ((~^(!wire63)) & $signed(wire64[(4'hd):(4'hd)]))));
  assign wire66 = $unsigned(wire62);
  assign wire67 = $signed(wire64[(4'hb):(3'h5)]);
  assign wire68 = $signed($signed($signed(wire63)));
  assign wire69 = wire59[(4'he):(3'h6)];
  assign wire70 = $unsigned((wire67[(4'h8):(3'h5)] << $unsigned((wire57[(1'h0):(1'h0)] * (|wire57)))));
  assign wire71 = wire69[(1'h1):(1'h1)];
  assign wire72 = {(&(!{$signed(wire64)}))};
  assign wire73 = $signed((!(!$unsigned(wire59))));
  assign wire74 = $signed({$signed(wire61), (!{(8'ha3)})});
  assign wire75 = $unsigned((wire72 ?
                      wire67[(1'h0):(1'h0)] : $unsigned(wire70[(3'h7):(2'h3)])));
  assign wire76 = {{(^$unsigned((wire72 == wire63))),
                          ($unsigned(wire70[(4'h8):(1'h0)]) >= $unsigned((wire74 == wire69)))}};
  assign wire77 = wire65;
  assign wire78 = wire75;
  assign wire79 = ($unsigned(wire74[(3'h7):(2'h2)]) == wire75[(3'h7):(1'h1)]);
  assign wire80 = {wire68[(4'hc):(3'h5)],
                      {$signed((wire61[(1'h0):(1'h0)] ?
                              (wire73 != wire61) : (~wire64)))}};
  assign wire81 = (~wire58);
  assign wire82 = ($unsigned({wire69[(4'hf):(3'h7)], wire59[(4'hb):(1'h1)]}) ?
                      (+((~$unsigned(wire78)) | wire79[(2'h2):(1'h1)])) : (~^($unsigned((-wire72)) ?
                          wire71 : (~^$unsigned(wire71)))));
endmodule